PK   }��XB�*h  ��    cirkitFile.json��%9r%�*B�_2��o�?�h��	ӳ� ݍ�ӝ�N�:�6*K-��ڗ�gZ㍈ʸ����_3FDug�(�2�i~h47�1�?����~�?�׻��?~����w�߿��p?�qx�S���?�}�|�/����ݟڿ՗����r_��|�6w��iо�CQN�Q%=�u�5�8�\���~��o8�!������	 GB`J��������z�ߓ����������P�꿰����'0��X��X��د
�����q��%2GıGĳG�+A�6�}���]bc�J�w���+?�4 |�B`*�@\�|����"��_��L�D�w�l�	�7:�|�|��q
�y��\M�����m�D���l����"�o�E 
��f�@|���(�~�-Q��]�D���l���n�����XU�o"FP�XP��5�:;��z!���3)I�f�
�ۅ������=)YB�����������,@�p5sCmO���s5sC��S��Ӏ�~����SH��@`j�^��=�@��Cҋ�x�x P< )7�\��{�p
�x��;�0L� ��/f��7�b"���� 7x��Q .�/|�N�R;���'5���VږNMx�ŝg����>x�x�Q�HD��3 ��a#�A��������xL �Bqf6� �>p3����N�����?��Q���_�Ѣ�"�;�L�n$�餗��}`gud�:���1b��3W��dkm����7~7�t��n-�P����F�("����8NS���5�lx)f2w���s�&��l���Z( $�,?Pa�8��x��M�X�E#�U#��n�{�N�{g�i*���;qÃf��ى�b�Y.�ܔe*����]ݳܸ�&Q�Ώ[�"NIrf΍�t��Jǭ�D�+�h$�x��L��t�n:�9^��qݞ�.�8���ˎ 3�>�L2w텉�d����忎-9n��K�`�y�D�_�a�@���-Q�W_�"���O�l��Ͼ�"6e�@|���(��q�D���l���;�"�w�E 
��d�@|�����w�E 
��d�@|߹q��}�>עH�8�E�����du'�n�냳.��X�uHh�����h�)Z�o��OUVV�V���8Fj�)�7d?��w��E��0��՝�՝(:�E�q���Dс,:}eueu'�d��$��$�;Qt �N�eY�eY݉�Yt-�/�s"Y| ��-�
�O�I#Q|m���D �a|��D�'�Qd�0��MX�LC�;��&�?a�!���w��f��@_��'�?a�!�����q"�f������& �>d�0���"�ma�!���������@���K�	�Y| ����֟0������>Sa�	�Y| ���q֟0�������NP�	�Y|˝���
�ˍ���
�Y|mﰰ����,>�w�����t�䰉��`_���ö�Wb��v�GG�T;.NBwT�q\���D�Q+ը®}�Cd5O�T�
c��^�v\���Si�qq6O�T�
c�h��j��Ih^�R�Z�/�;*7�n�՝(:z��qq�EG�T#v�J����Н(:z��Y�Q������j��wdu'�9�j�ŉD��\	F>�F8��fEҴH�I#Q|*�n�'�?a�"��@�������B�{
ݨ�)�B2j���,��n7�0_�5_a�C���vP���Ш�&<����� OD¤G߁:���O��,��ʙ�X&��� OD���I߁2��	��577/̽�Uz�
s/r����K߁*��	�/{iIzmI�����n�'b���K߁"���O�{��;P�w�<�	�'Y|��n�'�?a���	^M�VEs�ek��u�@���D�_���K����n���J��	�/�Z�U�����nVx�K�Ӌ{`$��o��UťҲ�kW��_x�L��g���O��O�{-�>ǌݬ0u��6�y�6�{ �=X�S]���
3?Y| ���
#�	2+}y;��&���1�%����,>Ƨ�=I���k��2q����/��&���[�d�焩�,>�w~���7K�ˋ�nP��۲{Lu	S7'L�d�0��{�D�'Z����݃��1�%�3Kzk���,a�儹��^��@�>�dND«n����걯�d�K�{9a�%���[���'̽d�0�v����ɓ,>��n�՟&O��@_�3QX��^��@_��QX��G�k�T
�Ox�J�k7l
�O����a|�nPa�I�.!}��0}�����Y| ����*�?a�!���d��'�?d�0�v������,>��n��_���@_�wXX��C�k7&__[�݅49l"c!�ץ��-�:~���?�O_����8z�\���*��ݐ�4wwy�����pl~y�������{^��ky�/��?���.��f�5;�����iy�4=`�0���L�������cڟ�nf���d�rq�UIuV&0n�![���Iͯ����z�mv!�rNzRbT9F��4�8&^a<��u�����qrC��
�j���T�2)��m��8���yJ���]��֘�0j��f5@�؃1�ѱ��vR��o����J������9X_G3���I�7�.h���
Q��]T�G�L��yK�曚7��Q�aİ�9��K�21�8Z=lk~����O��8fs�MSF�Y���� )�����_�-[��cs���z,ŕh�����_�<��T(>a�<���)���	��ͷ��o�]�I[��ڱ9~�*��͔k�\P�V�)�7l�}��Uf��+��!�j�-�2x��l�����!�T�)�XuF���U�?��Ft�[o'5��v�^��PTp�t&��|G�9�<z��mHͯ�=֜�b�q�ib�8�M���:����<���$e�O�j+��as�H����Xs�7�HJ��o���	�K�3$N�3����%����nk�I͙o�>A��_������v�M�ͷf�}�'�S��<��ƸS�oDV����;�Of� �=�ٵ$E��0����<m�(�7bjJ󍐚Ҝ��BGi���(�7�����4� s��\�d6\�c��V.�Ԟiy[�R{��m�H�ַ�K �g��V.�Ԟ������K�f�f� q�h�3��'��&��`�f.��|#�,�$�ʃFB�K4�$��N�0ŭ��|#�v�Ԣ�ҹ";�V� 5�0rw����)ͯ��̍�NA�T-���
�؃��Xǭ�����ۓ�%F7cx�}Q<e� i=oi��|�O�3DĈ�#�%�� O�:�y�	ưc��_;�4�&�ʐ��Ѷ ѵM"�M>Mj�|�������^M�������E�/AU�,��a�P��8��9$J��}'5����*�؄� �D�с�5�P=ؼ�wJ�S�o���|#��~�!$�p�0F�9�5�j����g������$Gi~��C�H��K�i�)��0�ѠQju��ik�#5��wR��}'5���)�h+�S�F�0�A�iH���u��\��od.)ͯ���|cܳ�)�b<26jVe�??�����͓�o�;��ƸS�o����5�m���9E@w��	��n�u�����|��Q�_��<B�&�Zb�F���Xe�k(��6�g��[kB��}'5���v�mD;I���H����������!o�u��~��|��S�op�h�����N �\�A�9�X�q�Ӹ�e(�7�w���;J��}���1�AM�-1N�n��#!�1�[5��F����z�I�7�=�c����O���L	�GM�s��(nUA��o-)�o���_�;F5�f�U!��l\��0;o�����s��)[�ܻ�E����Y���d�[3,���Q6�-r��L��!LE��䍞G���H�7���*	�V���M?]7����1Z�k��VWᴂ�Vґ�O%��R#Os.���x�{'5��|��X��qh�,ӤJ�m�i�&:.lͰ��ك���sb)ma�-�M��A����m�;��F�M�Q�� 	���݄_-~+��7�IH�7�>@���fk�U����"M�e�[�;��F�*�1��]���� C4_]��P'7m�	R����������������}�������%M��E%h����N�'���i�����lc}��vA� H���tZ��� ����!22��A������N���o��\���v�!rR:�R:��:�"!A�-}� ��j�"!A�-�� �Ok�B.R�k˹m!I��6-�I�s��떒�Ok�B�ļ7��o)I���/�ĨC��xȦ�����Ou2�.��q#�ǥ$�S=�&1?n����$}��$�Ǎ�������$�Ǎ���t��I
��7b~\J��~!)L����s(S	�#��C!"zt��ݵ��~��h?�BD���������P�G
�(Գ��ꀇ��r3Lz,<D����(솻�sN�����m���!z��։5�?�P�l3ѣ�yY��1��d��CtT����#xt��k�t��^��W21=��r����̞I��-)�B�d�&B���I�
���~�M��B��؛�i?b�b���C��z	9*&���)�"Wj��RH)�B�R�����$=�P$^B��I����C�y�2���C�b�
S�q!I�
�X4n���SE"�Z��=H���V̏KIj��JQ)+�I�K���q�l\JR��TLOO3�s� �� �9m�J`<H�b~\JR��Q*_`�r�N(�b�N7
ٸ��v������q'�Wy�$�]uN*O�������$r�N,��Ԯ��$�Wqb~\JR�JJ���b~\JR��H�X<������v5�&�x܋�U�$�+d�0��U����Ԯ:�$�ǽ���Ԯ��$�ǃ���Ԯ��$�ǃ��&��UԽY�0�K=ݟ !�`�.X���M#�R��+�`]����5DF���}H`�.Xa��.oF�*h�K���K��^/oL�*��X�V������>E��
]�b��E���,�h�V�U�]޼(.UP�=�B����FFq��z��`�w�75�K�k��k�	�C�0�.h��V��G��XW'��m����l���>h[�y��a_]�B��f��n�0�.h��V��G�}XX��m���G�}�X��mۋ�G�}�X��m�S�G�}Y��m��G�}XY��m���ga�/���m{���/���m{���/���m{���/���m{���/���m{���/���m{��/���m{+��/���m{D��/���m{];�����m�p-�ܳc�p\�����ǥ
�� �9.UP�=��O��{�׃��ԝ�]�z��Q��v��AnC��z���*�׃��TA���z�>��O��^r�N�.z��p}�q��z��p}"Q��q��z��p}"Q��q��z��p}"Q��K�k����|�u�����\]��O�A��n;Ѯh��'� VR�}�W���o+�j��=^�HUBv�⏪�>�����7����>4�h}"U	}��ъ?��P�.h��'� VR�}�X���o+��>�l�D��h��b%uۇ�uA{�>���+}x���D���T%��e]��O�A���vZ��ˎV�� V�n��.h��'� VR�}xY���o+��>������7���m^��V���/[��������T%��eG+��J��˺�]�O�+i�}xY��Dۇ��>�e]�B��n�>����VЊ�}��e�/�}�˺��>h�]5}t۩Z�/[A+��>��.���\�-��QB^f��.h��vR��`:�-��QB^f���uA}ж;���/[A+���e�/�}�˺��>h�a]t���.h��v�Y��ؑ}��Z%��e�/���mw���m�:�.ha��:m$봓��V�>����e�/���mw��m���.ha�D����e�/���mwL��m^�-�A�����>��Z胶���E��/���mw���m���.h��vk���e]�B��.�>��^�-�A�����>��Z胶���G��N��t�G^���2߇�uA}ж����/���mwF��m^�-�A����>��Z胶���E��/���mw���m^�-�A��T��.VR�=����?|�T?}��zR��J��s	T6���wC2�ܝ�"R��vP���D�x)ADJ��D�d�2^���#+62Vl�|���]+6󐧜'�'c���J��
0�q����ى$eW3$)���م<��9�I9�Q����`���{D���#����qrC��
�j���T�2)���8�B#����P��1�a�hv>�j�R�[c�c	vI�.�Z|�����G��ȭ:�����@�B��o�Ac�Q!�Q���*P��h���8ƈ"�2F�W7�0��:gTviT&��Ak���K��2�3
� �5(7M�k��.0��������b��a� =z�b ���A����@�B���es�v*��khuv�jtq����$e_/�Oڢ�!�A)�T.H�̔k�\�%�P��G��.�2;�Rq6BA��$,���L��(Rv�@��gT��_���1��0�0�'`!I�ł�A�E��|g�RfPq��cȣ7_G���%֜^j�q�Ym�8OO���:���I��k��j+�0f�	�2��tc�y���)�X<�sB�p���~��Ґ���t���$E�n�A��c�CT?�I��6�G�j�ٗy2>�Q���E�~�I��� �àlv
 �7��y����c�v�'Bf�"e��P�����k��}^M��O�)R�Y5E�>��H���$�2^�%d�Hbd에"���`Bf�$FƆ	�!�+&d�Hb�|���g�����1�0tǘ�L*�ɨ1��z3XO����G�%��Ay�� =/a�HMu�>��	�8E�>Cq�Ԣ�ҹ"!�V�h�ڞ�9k��dc(Rv����(��`�{Q�حI�XGBA���%i_bt3��[<�=B�L��L���	cD���g�\��G��JB�Cj�u�\������bA^����iqQ����Ю�sh��P2 $)2XvIʮ����Պ��U�"�FϠ*����0j���E�~&�"eW/$)�z�S�`���s���<:P�F*��)z�H��Eʾ^(R����BRn(�5cT�>Q��vH��a%Iٟ�)R�'j��]����W`ڍ����F.:h^�ls"��$)�z!I��Iʮ^����P�O-q~+v5�!ᯪׁ�'I�ςS���$e�^��ٽb�2JjVe��F?����,�;"Iٷ��}{�H������ۂj��~��^�g5Nc�S�Ļ$)�~�"e��R���e�L~�1b[WaF�b�6�5�\�W�+I
aՄ eW/$)��g��R�襒kYR��Ck},zȄx�$e>�Hٟ�(R�yc���XU�	g5�*�yPq�.�a��4x#E�~��"e?�K�������d�z�0�l�Ơ|A���L�$$)�+8)�z!Iٷ�<�qD�7��Ƃ.<%tZ5�����H��$I!�k�*PRv��P�#F����C���nA��8���jE��<mt��i�L[ô٫<�;o�|@�N�(R�WB�A'�}h�<媆05@*�7z-�O����GS+��Z��Dϐ4�7�@������Iʾ�V8-����}�m��
������U�I�����5Uǡ�N�*)���Q��,�@�HR�sA1%��RZ-@[g���̃6���#�Iʾ^L�Q��Ud6���݄�?�IC��?��},4+j��eq�C�"�C��Lm�5������1S�q	��P
:�0f��%?ur����<��'1w_>���e�R�}���b�}��y���|IӠ}Q	�0	���S�����r�P!����~��9���@J�C��"!A�4w� �O�"!A���-�HH�>��� �O+�"�����"!A�T	 �HH�>U� �*d\��זs�b~���$�P�!�I�w��󖒤JDd0��os�R��C�&1bN\J�~(���$�Ǎ����
~d0���r��7b~\JR�9R��7b~\JR��P��7b~\JR�O��7b~� �xľ�%� $��C!"Dɡ		��P��SH!�w�ԃY��\�DR��.�@)D�HH%�BD$$��C!"�ل��E�ym9�-�	�*&1�M�|P1��nB惊I�{2TLb�����b������'d>��ļ8!�A�$��	�j`)��	�*&��[. �����'d>����8!�A�$��	�*&1?N�|P1��qB惊ȈKe>$s(V̏KIj���a��V̏KIj���a��V̏KIj�\�a��V̏KIj�*�a��V̏KIj���a��N̏KIj�Ɗa��N̏KIj���a�ˉ�%������R��m�b������R���b������R��mybK?b~܋�q)I�v61Lb~܋�q)I�601Lr��r˛b~܋�q)I��&1Lb~܋�q)I� 1Lb~<��q)I�V1Lb~<���k����Bݛuy��ԇ�`�B����[�^$-UP�=�B��nqs��TA���
]���m��R��+t�����^Ɋh�V��.z]\"+��X�V�Q��uq���z`�.X����Xi��z��`�w��c��
�V�U�-n���*��X��V܇�a\]�B�����n;��N���>��0�.h��Vk�G�}�W��m����>�Z胶����m�-�A��0��m&�-�A��b��m6�-�A�����mF�-�A�����mV�-�A����YX��˺��>h�^�>���˺��>h۞�>��"�iI�/3}x���˺��>h��>���˺��>h�^�>���˺��>h۞�>���˺��>h���>���˺��>h��>���˺��>h�^�>���˺���h��{\�����ǥ
�� �9.UP�=��O��{�׃������^{`=\�x\��^{`=\�H��E�yu�Y���z�>�TA���z�>�����^��.�.z��p}�q��z��p}"Q��q��z��p}"QI�q��z��p}"5��C��V�Qc�>������7���m'�Շw���A��n�P�.h��'� VR�}�W���o+��>�����7���m������J���x}�b%uۇ�uA{�>�����Cɺ�=^�x�XI���e]��O�A���B^������J�/��x}�b%u�iI�/;Z�w�XI���e]��O�A��n��.h��'� VR�}xY���o+��>������7���m^������J�/��x}�b%uۇ�u�O�}x���˺��>h��(}tۇ�uA}ж;^��/���mw���m�j�N�}x����l^�-�A����>��Z胶݁�G�}xY��m�˩�n��.h��v'U���e]�B��n�>���˺��>h�a]t���.h��v�Y���e]�B��ζ>���˺��>h��s}tۇ�uA}ж;����N�N[���2ׇ��>��Z胶�i�G�}xY��m����n��.h��v�d���e]�B���>���˺��>h۝�]t���.h��vwi���e]�B���>���˺��>h�]�}tۇ�uA}ж;q��/���mw���m�S>:�ч��>����e]�B���>���˺��>h۝�}tۇ�uA}ж����/���mwxw�m��˺��>h�]�}tۇ�uA}ж;���/�hh�������˝���UG��K��qUEW������r���R��'"ŋH	"R���$"%�X����X/Ș/��/�0�X0Ș0��0�1�X���b#�e���Z���<�<�<�\gUR�U�	��f����N$)��!I�U��.��IO�A�*�蕝Ǆ侮�#�������Ȍ��\TU+7F�2�I��ؔ���Q���ȅ�m�Y�F��iV����0K��XHRv���k�uT%�=�Fn�)����f ��}����
Q��]T��G�L�ƙ0F)�12��Q�a�8�9��K�21�8Z=��h_�.�	��P y�A�iʨ]��Pu�a ����$e��ѣ��z,ŕh��],󘳶sP���\c@��ST��h ,$)�z�~��JA��rAd�<X;�/!�"e�;j�uA�١����
�$a)��g�wD���rH=��Ug�|F���7�)�}8I�.t�E(�8�;�g�2��#�C�!�:��],���R���js�yzr贬שd@��HR�gX[|xV�X�G�1CN��k�3e��H���Q�: ��=��3����%�����`/$)2Xv#���ӎ��)?L"N�y?�P�ξ̓�)ƈ"e�^(R�cL��}�e�S 8�ٵ�S��0����<2C)���"e��P���e�XS���j��}ZM��Ϫ)R�I5E�>�&Y����X/!3D#c���I��2C$126L����X1!3D#�e�x?3d�d͌1�;�DfR�OF�9L֛�zJf�$e?/��8ʃ�(�y	�Fj���i�H��)R��Ӧ��	�h�JE{����YS4%C�����-E1S��#�� ��nE�H��:"��],I�����x��y��0e�f���L#����8CD��D?b|VZRӬc��`�H�$e�4�H��re�-�v�C��!I����`HRv�K5�ήV$|�*�0zU�V�QC%d�(R�3�)�z!I��˜*�؄��L�с�5�P��L�Eʾ^(R��B��Ue?��rC	8�����}�CҤ+I��LM��?QS���e(6����n�=��4r�A���f�a�&I��Iʮ^HRv�2�m��|jaЈ�[�#�9	U��,8I�~�"eW/$)���-��Þ�Q�P�*S��5����g	�Iʾ�P���Eʾ����T��S�R>�q�0�*%�%I���)�~�"eW/�e��C�ۺ
3j�q��䊿�dXIR�&)�z!Iٟ��8ۈf�jE/�\˒�Z�c�C&Ļ$)��E��|D������ƪ�N8�!wP�̃�st�㔧��)R���)��^��]�D����&��S�g{7�r����g'!I�_��H��Iʾ��q�#�a6�5t�)�Ӫi�t�FB}$I
�^� �P�B����j1j�6��B@���v���av�V�(R��i�S�Ncg���^�	'��x[��uB�@����:���Cc�)W5���R����h	|�$e>�Zy��
='z���G��"����'PV�HR�m��i����x��Kn�VH��\����_HR��(�e���:m�p�TI�����Dg�B�@����)i08���j�:�g�	n.��^HR��b����
��"�)U%�&t�Nr������c�XQ�5-�jy��Efjˬ	��$e?��꘍K�̀R�A�1��.�i���\�$�9��|����_�������8�������Ǐ��ǻ��:�}�t��~�����oV�&bU�3�϶���A��4���\�Q�Z�����N�]����ۡX���
t����a*����*�	�
��8����l���]��σ�e��9�>�8��`y "��l ��_��`ڠ�\ �y� Z����@s�z�)��r@��*�5V�R�4'���+W,�C#	[^Up�m��-������o�OL���'�LEH�?�0m/���?�1g� �'�L�s�}�:��%䢟���~Qgv���~�o+�>\2/��å�W��ַ�پ�f�^�ix��-s����I~�|�~f
kJ�&�v�7vf�ޕ	���,��A����-)QC=~Ґ�$	�� S�Dd�Ɖڜ6NĮ]����E�\����E�	��Zj��ϛ����U\��I�з�5]�<l �<>�C�1���@�".��H�	\8���X�v.����͂�2�����jw�����p#a8�b����e�ʤ��i㫙�W�5*��������L�?�u�I�髛�9Sm�-O���io��ދk7�"W��z���D 6��LVw����>E��J�:��S�V�4���  �@;����9! �3�1�{؞�=%� ��:�wxm���fD6og�a~lƌ
�9)�Etx�:E]�0̕
�d�D&� ���,+��Ģ��~k�8���I�c� ��K7�a��u��/��Ҕ��Y9m�/+�-Sfzei�a͚��җ���������_z������� v�e1�N'\��۳y/�nJ���I��E�-|;��ܕ�c�0�>�����ZD������j�7��n1\w��4��9�.\�s� Ѳ��ǆ\��'^��K����:��4������ս��_���c��X�h$��]};� ^~��jh�xZ�%H����G@]�<�*���ކ�;i�	�f�NZ{ٚV����X*s�] ��n#[�ήk�Lt]�ܠ�(�[�'�$�4�g���.8]�:|О�e>,���+{T���g�2I�U�Ç�~��f-m>�ya&C����"`��3���*�"�r��t~*����Τr��V�_Ac�����M��u��b0��}0W��O�*>�8��[��W2�~؟D �VGC.���b�����UUݴ�"Z��-�}8����B����E?�m<��U1��|ܖd��fXή�aNq�_������'�b%&LG��0�"% �JV�
|�L��^�b�7_�G�`�1�~W���G�~����xk�<^ݧ�?`�����Ɓ�t	<���1�,0�a�]r3�e���uR�;F�8�F�=�}���jv�s[�嗩1�R���s�R
��w�1���d4���jQ��]�=z������z�d�������>�[��O���j�A���r���"�K�N�ސ~����HZ?����������9�[ ����+���倯mB� S�K�*D�ep�ot�����M�p���!,m%H���Q���]�`�<^�w���"_{Z��7��W��WMY��k=���B�oc�VƔ����
����4�ӫ�oP#�
[�1���4�ӫ�_��m��u8[�1}��*���46zzQb��nc����U�7�D�uǿ�8[���lH܆X`�7�>K�p0u��w����op�\]��㷛K��t���ߴ.�	.���Zeҁ;�Ep0Y��B8$B�o���"џ�߂�L��q���r�l��Ϊf�}�'�N��0�A��#���E@p���m�����z*�1�>�v���E��K�r\��x�I��㸩B���/��CE�F���\+��D��W7\��_���M�Z^WE���W��5k�`{�[Y�k;2NZ���z����z�.�D�k�9�\�_�s'2�L[o'��?s�+�?	�N鳸���~_��ʹ;��K8�+}}sU���.����������oo��>�wqk�$B<teu[�9�v�3��ߟy�u
Bm��t�7�������p��0��!"[��D�"�ᘔ˃�D�4��^��.�n���H��K�`��E�ZԦ�ʸ�jhb@��ͺ�݀J�[4���'�I��J��J����T�輽�1��s�Wm}m�_.�,��cZa�e�R�$��j>�FO��h��zA�%����CZa�e�8�S?D��x:{9O�|�Km/O{~	No���2=�Ne=���N/�i��z�����e�DK��<��˧���]p�,�c��+�<-p��*�_���(�ρ8��� 1�waL}-���޹W����k"�$�1	 "���S�y"�y��-�-)��f���4!�}IG����|0}S/ޞb33�ݒG7?�5W�\��=���d]%>\�UW�5?+�to_�B(����>��?����H�y��l�x!(�'�S�񘆺{�;7B�=a���K�ƅ=ň�8�WK恸P̕����X�U>��A	7e��E�K12>�>��پ���%�2��E��uA��.o7���/:Dż���o@�A{y{�*�ܶ��\�6�ˋ9�1O� �E�����7��tżA{�_�1� �+^Q�5��܂��xW�_�Wlkg� �'�t���K%x���՗f|��XR�����Ʉ�ͮ��Ĺl<{��T��ǕAhE��R��ri�!O9O*O�(�Y�Tg`����g���\��2Qw��Z�ʥCv�hv!��9�I9�Q����`�b9W��B�&��"L!��2\��qrC��
�j���T�2)��ٔ�ٔN=����ݕ�n �E��`�~%(;D���e�F�5ì`픱�8{妒U�V&�9���5�+ �
����~��L�X���� )$n}��Z���1I��Y��Z�D��*�V��(�e��+�xQ?qm���8ڬ��rC*�STc��q��7W<�A!܂�=#�X~]z����0��f�l�c)�D3����! ��~vB�&���N�:�ɢ�r6{���Dg�m��]� 	�̈�m�>+�!���I�־�	H��Yk��ܾ�iQ��[̵s�^w@�u�˚�t���n��Jsi�_�n-��XGU"�4uT�B>���`���y��Yp���1���c4�rUC��� �L��y�Iĕ{�H �&�kڑ�CĵdM�H��Q!j�D���x�0sM2�B����
�� �%�Vv�1�I��I���yN5�ߊ$��!6��V��`�)D>�މ���1E6^b~C7?!��EE@\�TD.+�^���\V����۽����=�e�rgܜ�nF�g�eS�ܥ��7���({�Iw�I~K�����L��஋�h�K:D@p�.��C^@��K|�*�p ��ʜ&���X8��9��{������J�R�UO&	�`��<e�2L}��\�%�/�ÈY�	�'��~#�*wt�a'U�"V�-U���֐KU�rk�E>d��#�2_0o�8���&<)]YA]�\���6�	��R0�K�m`��R�8�a���Al.�F�lŪ-��I���k�bG�0YՊ�{c7�	9�@�;���Kaoo_�5T7���*���ʫ�V�Sx��1Ch�c��Z������[��)hB��W��:�v���{l��2n*]�A�;7OnK����Bb�3&�������*��~�$��<���ێ_u�#	j����q��C���W�ɠ^`h�n>�5W�%G�0������%�9>�fJ��۝c�S�(��qr+X�Nv�<�M(��v�j�E�Ջ0���;�����p��e4"X��ڹA�����r�E��7��J��OyH]�g7 [=]Z0d�8�M�Z�����zT�էV���0�Ȥ�U3�$H�3����m�G��o
�8�F~�đ7�8���n�H3��:ܘp�%�wy��Y<���M�[K.�5�^T��?�#�Xx���B
�BX0���NHL(V��T���f&��;�u	�3ǅ"u���i7��7�h�]��Խ��4w����P\Aǋ)�ד����܅#��W^?�İ��Y��2�en�8�ũ[�
��{��L�����s��>e�~�������w?~��w����������/��~�8���O���%M��W%��쨒��:�|�|.m������6�$�p�x����8�8��UVEe���6�D���)�ה]���)��x-�"bt|My���"sc�`�hq[Dc�llm�e�`�8�|�.O��J�^�����  �t�#[��K>/
n�/㔢�����:p� �[�2t[.�/A��o˗qJ&�qx[#�m�2N�X>ok�-_�)��!�m�����8����!�^��{��8�)�ql� &-�I`��r��E�(�9e�Ɍ�t^J����+nˁR3j�~1�,�9v��B"7���܉��h�9���#3{�"�Y�������_J��u���ȴ��L���u�+�����#h�d~5�t�ܳ&WDZ�=���$M�8V�?sUt3�B�����0e3�B/�X8Pf��a����O[�
k+|��`�x̰\��9�o&\����<�%m��m�w��R$�V*�
kŭ3�H�d	�?\B\yK�ύ�7S9TXl��ʹ���F:��L�Pa�=�N���c�;�.K���Fw�@TX�a�Y�o��� �ە)�[ǳ�sK����SE�4���"�\����+�!�	(+�!f^ò=4<ȸ�Ŝ��J��=�u)�Kn�J�_��dBD)0%�e���V`�����  �t���_p�x\	���R�@>�-'6�e��=�kE$7��V�=��t�u)0%��)��:������|�'���2�@z�/C�y?Η�8�s��!��2�@<Η�8�.|�C���e ʗ�8�)_��|�C���e� �O�2��?��h��X�x���;��Iym?3S��v!Iy�����'���.ȵ㇨�~��4�p���%�����]�ev�
��
[����	��"9V�V�,>Ƈ�������d�0>����'����(��(�?Y| �O�%a�%a���a|�.�/�O�k���Ѷ4]F�[����)�8g�E�ʐ�u(��4B�F�J��u(MN��4�V�-�CiF"������et(MK�.B(�Cij"����K�P��#i����yJ3a�����]�&)�W&�,MS��� �ili�"����*�:��)�A��)�2:��)�A���	Q�2:��)���PQ�2:��)��~*iJ�a� ��m��֡4OF���5iJ�a� ��m��֡4OF����Y��v��eT�0 L=�j��	�;Pv\������<����-�̫R�LḼU��;Xe�(��V'�3P7��xK�etJè�V��I��=1��(��@i�qy"���w�4�ZO.�?2m�֪�O߁Ұ��D�'��@i��d�p\���d�(#����q\���d�(���l�^xE����0�#�a7�ѡ8g�Ex�4��2:�f&����� p�뱮r?R)v�@�J�z���E�J����c� �)�j@���˲�]�&.���� PF���E�±��P��,^�F�lG��n(�RiN#��H�Wg��Ӏ0�#eeTHsz����Gᑲ���*�]�_���<��ʘ�4�Fx����2:��8��T�� PF�ҤF�*���P��,^���i��,��X��Ԡ� P�J�)��ei�#�p�MP�j Ī�Y�A�T��Xi�c��q��4�v����9�ṝ[nu�4�Ҕ�J/�#i��*i�לIs�%�;�v�UҔ�.�E\Ĝ���
`����f@�Aa�oCZ�;���4!Z�j@�Y�Ua� ��]]"�CiʳDx1_X9�2*�f@Vz�G!H#lW���ISa� ��]w#�Ý�,��%
��\HS'My��4�v���w0+ل�
`��wڈo��k#�q�4�q�G!H#lHI�Pz�G!� ��NY���.,i�Jsa� ����%�Ci�#���;Ȥu(Mj��4�v���4�F���o�:�^�F�۽u�:�f1�Aa�sOZ��7�Aa�/PZ�ҴE!H#lwJ�P�� �c�i���-^��#i��IiJ�a� ��ݏ)�Ci�"����=�u(�S��4�v/���4OF�۝��:��)�Aa�v{�W�֛��˨�+`�<~���?�O_����8z�\���*��ݐ�4w��9�`�ō��/n�=��2�/n?�~qC�������_��}���&��7`��r-�&\��
�k���C�"p-�p-Ѱ}!�͆%�y�SΓʓ1��qV%�Y���i�l��l@j��R���B����Ĩr�^�i0qL(��~R������8���E�P�rct*C��iӺMi�M��?��~��5f5�ȧYP*vb��`t,�n���~����bU��!��`�S�±��h�|?������Q!�Q���*P�h���8o��~[��W7�0��9gTviT&��Ak�����x��nb(�C7נ�4eԟ�j���0�B�z?����G�h"�T�ۛ0��pm�c)�D3l���~��󘳶sP�������c��F'� ��Oj���'m�t0�����\0�7S��rA����߲���VT���艇P�#Fz�r��}޴J���C���R����3����)L!��E7�Oj��~�|��PTpu&��~G�9�<z��H�7�kNa@�1�8��1W��&���z�J� ����~k��u��f5��ο9a(Qft_n�9���'����=jl��T����A�!{5A	>�l��R{��7�oR���ˎ��)?�n��Lђk�ٗy2>�M�S�o�?��V�Ei�ń��fv
 ���]�s�Y�C�1i;��f6��~+���
�)���"���[<��~�R�o�@J�-Hi��I��6@�nf#H�6��� 	�Z�f6�$�k���� �%nf#Hؾ�k�[�k&kf�&\1�0�J~2j�a���og#H��JAު<hdӀD��A#��M�4S܌F)�q�M-�)�+R��j�
�j�	}gM��� J�������)(��E�U�H;�"��9��o�?i_bt3F�޷h�#�P& �	����I���8CD�H�=�y]����c��`��(�����1�� �A2�l���E���sh"�l�qR{��7 ����_M���鋫�E�/�#AUd9��a�P7�A��[�(J�����o�N��
lB6�����@�]��Nm��?��V�)��Oi��d?��rC	8�����}�C�;�8R����~k�����Pl�I�]]w��hdS�F���6�����~�����'����R���#�$Ŏ��4$�U�:lfCI�����'���lq��0��퇚U�����nt�8�i���[�Oi�5���[�/8��c[�*8N����i��|���������������G(ӄ�N���U�QΌs%W��v6��~3Nh��R�-�o��F4�T+���Z^����Z��f�Gj���)��?����֚�*:���Ѳ�eT���e�<�����~+Hi�������ޏ�j�m5kp�tcP� �	Y�yތ�I����'���<�qD�2����N4%t'5���ç�Y�Ej���Mh��Oh��j1~�6��B@��V�
j��av�l�P�o�F�lR��V�l�*O8����:�Rnο��[�Q٠��-`n�1媆05@*�7z�&�#����S+f�Z���7i���Ԧs�~��>l�F��o�_�Ӣe[�G�>��fR��=͹�����~K�i.cE�Zǡ��L�*)�լQ��,��9���o�bJN����Զ�7��m��h�9���[�7qp`G���5���w~���Lr�^�!��z� �T���i���PȤ�-r+[f�����o�R�q	���=��0���%?ur�&� �x����������;�����R���߼k�!�_��U���y��p�v�I;��]P�ۓ����銀�񸧳�N�@k ��i-�Ivka��ោR�sX؈R�hD)j��P���Pʆ�P�|.!��5�TҜ5����5�Ԫ���P\r�%B5�YJ��YJ��YJ��YJE�YJ	��smo"���6�����������>a��ܾ�g(g(+��9!�ր�#_uJry�!!+�ng�t�jCJp�!%���FB�i]9���jCJ�c]��$��� ��ՆZ��F�[mH!bg_�9�O�s>����D@ ����� ���o �����$D��`��C���~i��������N��9^~����\<��U	���O����S�����r��ۅ-o�X�}���a*����
8 ���N��:���m5�6�џN,|���\���1VYb&&�4��1�L|������]�D�D{Mg��{:�,|׿Sj�=|���{z��w���M֗�v/=�e"��UP�L\��B^�i�Dȳ�v} ��i�K�l��u-{�x��EL�y��zȜ���5�l����K]�C���C_^�@��ͱ����K���{���5K��Q��Q^ލ�Dx5����y�����V_#h�P�bNb9�2�j�Dxy�
K��
�Mp�h}��
�˳�y``EC�0
�9�X��*K��&���7I����<"�Y;��%f$�V0�.\MBP1�ؼ�b2̐m���w�zZq��M�Y���%Bnh�u�y��iA���dWhϡj��o����a�b��v����q��v��
&��X.Tߙ5��bbMкmB]ꉛ��]S���e3����u�8���eE,�ֵ�Bυ�;���n9^��v�L��H��:ߗ��_�J���T��������y�m����C�h����_��_���I��W��Wy�+��+�����_�*<�*,�}�O��wO�`����`�:x���S`��$�,e�'%����Sܲ��}n�>�$ӭ�|��dv���,��'�إZ쓪�R��Ɉ�Ҋ�ϯ[y�S�����{v�=��;��'�f�������'U�U?��-�	?@+}����SvO�ܲ�{j�V\���`E�ϟ�Y?����'}>��n�}7O}��@�6|���3���������?~i���Z��&U���|UI�Ne���8�>ݙ��u�SŀU�����ׯmm�����;:��9�����uh���)�Wn՜�*Sj��d2���Iv���|����e�f���A{��;g��?��ￜ�J�(����;�s���3|iU0:���?�P�|����?�����Z4����Բg��?��߾�o��?����'|a8}�?}��y�����?��>�7���y��Ǌ�������?����?����O����/��ç��a���}�߂����X~��p����'(�I��/?�*~��ȂN��(�{�R�2:C���Y�n��w(��d��Y���<iUk���΢���w��w�F�����W��w?��e�4>"�ѿ���#J�{4�����}}��(���ȴ}�d}83�߽��3;�h|tP~�`>=��Ã�A�1WLS�&)>
��7�+��GA�Ѱӵ݃�d�|��̣�G�@���y�q����Tl��'�b��s�����?IW��8d�<�$�+
\{.ه�R|�aX��ck��|�_S˚�5=�>�2n��]\{�a�>��BWX���/�}�k����ߝ������_~�>~��Q����ŉ���m�o�u��4��?}��W�i����?�{q䃱�h�G(=}1��}{�RQc�*C;����0�`g3��7i�ѥ��>����}���`�Mx�t3�q�Cv�~f�]�^�g|| 9��|������O��}��\��")�~��7���;������%��1�C0�}��]̏�s�d~z��m����ڬ���l%?>��U>�����`�!���� ��l������RlM�Q��� l����=�E���,��i@rA����a �bJ!��Ѽe�#�̴?��u���n�?�4}�~��a&9�K������d>a�{aÆ�����fϤ�8k��4�iD����$"�f��`0�6q�U�ɤ�ϳD�hR���fR�&��3�taL)u1&�Ng�19g���p:�Z�K��K1��OF���S��NI�<�8�9����=U͜��f]����vH��i�c��v���Y�IKK��پy!9C
io^��HG"��)����h.#����[d$o@ܙ�g������	$��֜�<<�Rʋ([ʖ�g���Cg���������G��C_Ǵa�:����{1�m�.G�����?�O������Z��E�nZ	����}����U���S_�����CS�����G�<�u���M������e�\|��?�z�W�0�կ�Oӏ��.�}���{����/���[�.���%��ql��*�`�v5*��*�ٹ8��Ӳ�3]Hk������d�W�K��o���x'c��y0>ĨS4:��?������_3�qY�ͥ��H\��/����E�����-a�cp������"��#lZ|���l�/�vA�����%b�Ql4g�@�@�2��ɪ��_�!�aD�N�aާ|�:0k�6�g�]�t,"�!��p�3�!Kˉ��L�O��ǈ�=��̨u�2��'��R�4wg�_���1�=<�K��a����\�/4�`�ˢ�m.�~@�c[����O$�J���*;+ʅ�*�-�|��f�� N�w��=S鈁uD7�N���Qy�y��t<}!�*%�+KrV���Y��Y'��B���<�Hx���\L��T�(3"�$�r`/iD��K�=E�����o.o�~���o��U^�P�z;���󯱃�IG����
h/�Eu��(����\�x.\y�G�s�.d����
�]ڨ�h�cHO���s�����-��3*.��rHG����M��.�+�>�)��n��g����e����>�H��f���雿%�I���s+���s:\����ؿ��T���N���b��n����z���(�\��î��*K8��S�,�Qa��C�w�l������C�~�Ӵ�<mRq��Be��^����a�I�מ{tc	v�{ڔ�TPs�9��kh��1�|�й�g�n���+��������W�{�d ��]lً��ZYn���疣����
V�[����V�����ן[~E��-���s�2I��L��*�	H��C��Y��L۲gZ��ů�C���%�D�E�r�9��#�e����e���o��e��<`�1�66c��`,>�ƥt�>wJ�R�@��;<�篚�㮎���/�ȅV��:�`|�1�l3��i����b�K�H6~Z�z������/�*X|����k�=؀��m��COR_M�M�b���B�������)��w����I�Q���%(���Vk�������Ў6�*?�*tX����=���s{;� _����О���,�#�/6B��I3�4
�6����9�{F�����7�{2I�:|�/�.����p�7nUZ�	�~d�h�t!���������?�����ֿ|���2#D����dU�+3��s�d����e�V����>����ե��ߵ��ғ�?��k���$~���Αۛ��������A��}F��:�\�N+B�{
�~,�jV��K�k������{����������7����?������vH�C�ڴ-��R2��'5���i;U�h ~V�5�<�Pk,@,��\PM���ᐓS�bs������C�>2��þ�}��#� '�a̹�8�M�Ӻ�_��7�����^ukЌ�=��S�\3"�RO<��a{�ї�j_	�_��7C�2$g^��S;�Rke�)v�H����o�B�s��Zr~*���r^��������_E�����o��Я�?vJކ��ن0"޲�V�>@Q�����f�3�4#)�J����b�۶�v2�o�5��`�LHs.��`����D���Q�8�����26d�~'�v��V�u>���!��� <7���j�Z5"�R��Y�m�3F1�F`>$L���\ƚ�����"M�*)6f5j�D-�@,UNЦ��}@)�v3>�a�_~3��\��q1%���Ngi��Y�<h܌s��F?�a���_+��ÿ_6��S��+կć<L;��K�(�88���X�*JUɻI��A�ϑ\��5\���G7����hnL&}��_��Ct���?㑏�>����.D���0@#E�ִR��p/A�+�t���z������r�'�W�^c�o&�K4y�O���K�c6.�l̀�=�v�ƨ|u�OC�ܴ�-|Ų���O����E���!X֩�Ye�s�lni�`Tyt--]��K�I5��$X���-_�E^{�����
�^�p��A��ˎ��ѪTki�Z�!����Z�2� 6-Ol���X^����X�m��/�K����"���Cyx;G�G�?�:wq�n�!ک�߲��b�]~�\�[b��yv���}(���1f,S����k�>��;t�0���ǌ�Ӧ�����`�JE{0��;���|õI��G������c{���/�z�Ϩ�w�Gz��N���0\����q���&#!����v���S4�?m'&�ɞv���e���x�8���ӯ~�"���/��O����d��-������}��o�����������������?~��w��Wkל�;{�W?M+�~���z�ߓ������������?�D���.Z��OE����qO��{?�?|����?_~�����������0�c�ůOy��O��M�����;���tG{���c�k^<������D�9H���D�_���o���O�_z�{���U�Gǿ]��|dc����ϹKCY7 ����yi�R�`M��=Ȁ�	k���k�j�-�����ko%��y�6Va�7��4���
J߶��EC~�����=����y���̪i�s��{���-�n�Ef����c�a;Z�q�h�M?�#;�'�b?���b�o�����y$���=&��O��C��,��:�H(��5��fWz�I��������C?8����|����/�˴/���}>Uڋ�1�;����}y�Q�j ��1�q� �)�4nʁ�q�NG����9��S HZ@�B� �H|X�N�@���s�i`����I!U��߰�B
ɰe���Ōn�|��ϝ���4.Y!���{_Џ8Y?�^ʏ�~d�A��@r#��^/��w6���/d�"qXԯhCc��^��0�|1RكU
�JC����^����2���V�50��r��k��dT	O���4���������_�E�ח�_��L(m}�7�P�,��"P�A׷-0�|���Xx�n�u���rq��yﳗ�6�k_~&z����>�B5�2,���s2����1�r}���+2i��&
�!��_�Ȏ�U�|�U�
[��7s�RY��5j���
�Y�kY���^�PJNM�K�؁P���NW	��s�j[��=�2��V�s	�����s��U�P�ˬ34�{+W2����_���`�]��-���.;{�!pȐ�E�]��'ePPR�!�c���~�(�]1�Z�A��L'�nX�_�5yW_��ҳ1?��������t��f$����;ؕ�֟`<N�ם��W�t�W�n�� ���#k�Nv�p��88�Dy�K�yc�@��L������v�с��U�c�aU�iݠRb�bX�6��ҵk�.U��������3�Oij'bz��޼g�]����7����2D�������ƍ��F����; ꘭���f�L7��q����4EǊ-�iã�ؽ|����'[u���Fe�!Ƙy���u�*�6كA/�4��e9p�rؖe�:p˚�n�d����,BV!��������`Q]��fΨ�V0?�������p���+UDh`�<��r�LW�e��ա9��j�#�eR,�yE�3
� "��F+��)��Y�+g�6����,~qk8;�W=fR�:4q&c���u��ȡ�=�^�q�iNu�7ԒV�#K�-Nn3J��׮81 j� �j�-�� ���2��*��y�b�.lb�7��cZ�V�!�����T����l1��,Tj2��� ��d���/;�� j{.@���ddeFX"�l��-�EH�N\�"B�K:t{�"Du4h��@��D#�(B�Z&����!ԴL�ha�: ۟Ο^g����z'>{F!��55+5�EZ6!zK���U�h�T�2�}{�*��	@�Q㋼�����w≭�:���@O�`�f��@��_�Z;4�Tq|�J�+��E��2���6�u����Ho�^!��`L�
�q�z5l�&TC��*hX�L"ԍ��6�I�C��D�;W��P�p��KjQ]�(���(4N�g*Qa�c����R!�Q`�LW�c�y�
B�C7�����<���n��>%���v������׸�����4�ӯ�=��vx�1mN_���{�|����_PK   �{�X�����   �!  /   images/00133a18-aa29-496d-ad09-d18fc42e20cb.pngmyg@SM�v�&(��EE@B�*�(��ޫ�ޤ�h#M:�""��  ���^����N�?�������svgg�yfvgO4L[����USU��.��GW(�����#w�jAA�
��S[
�M�j���I�KӎlA �5E�AP��T�;����ʆ�#8�x%�A�w�Q���6�r�+/��K�^)�C#����¸T͠ד���|�3�<,��,N!K�CW�'����ǣ#��v���-�嬆J�X攬����6ϭ�n�~N�-'�"N�T���c_0��	����|�����E���}�{lW�P�e���Ѥj��K�x�mĭ۷���t��7�}��(�#����� �!\58�8u�/��'.�L8�X�O��
r�g���,�C�!?���t�(���͉@^�7v���xA�(]��l,0ɰ�d�ge�b<\�$V'p\�������Ok(������[��4^I��G��|p�n����g��UV2�3a�8��DD
�J�M�?dt����N�%�L����j�(5�QM�>^��\T'�����&-�b!�MR�j}��^��Sc#��t	?�	�d����t8Y�^Ⓦw�B�ݭ<lְ�30}@��\���>~ʘ��Ӊs�CNT�K���>�y�^v�����Mb�0K�
�&���|�j��s��9<h��"/Z\�dOs���Z=�FҴ>���iV��
k̍�˝�b���Ff�䜅�TX����P��:ϫ}p7�����Ժ�<A^�i�@�/A��HՓ�"�������� ����q���]�QS�w����Ȍ�	�/�[�3�״�����a͹`3�$W�ayP��i�vwL?�d�����R�e]�Zʻ�v�⩍�7�_�G�G-N�c~9�6KYpD��U�4�_�]��g�+��.�D�,6��Ȩ���'yE�<%�"4���_��/h�-;��:v��ctR^��cUJ8��tBc)�� �Y�h�dǙ8���`{�Q/���se�c��~�a���B#��=����x-����$��Evz���j���S��@Ye?'T0��>cd}�s�dl�c� �e3MC�h�v?'�\��)&-m~�\�&�eģA&�i(��RG-a���_քck�(I�^
���4,��@�XǾ��O�oia�-	�zy�����*%S"�mn�&Z^��+���H�v���`'W��|��0AG�܇����#�2|r��K�.9�����Xp����'��դ��ז��>WL��B��Z����z�w�>�����-�u.�6�`KT��\�-(<*2��r�����5q�vR����pxd8�#=?T�`�c��'R�K��՚#�(�=z�%HjĚQ�J�cV��ޅ1{z�GIԓ-�*��zx;\K9S�ZE&4ť	�m���#R��o����^߈㓧�W'����uА��+R��v]D�w��[�@���^��[�%!��W���DKK{?E���V
J�eq �ah"6 D���)�j�ܖyK��Oܺ��Z�`F���&O$�W���a7]i��o��VVF'aV? �1H�N���8<�GoD�S����T�ƙ���]���k�|Nzf�}��|��1?j$�C>�æ�����mwt`�2y���3���۳�����m'l�����?M��v�Za][A�s�N����d<��<?/��C�{�&fdm�����	������5��>�L6�l��=���rR�'�9��sS��'���h(&8�8�r�V���1Ԝ��&���:��Ǔk��IGc���0+B���z_2����MR�	n�AZ|h����e+Q��V��P@@ �� N������F�4�����:G��<�?;;�ܺu��+**jdyc��tg�b�s�t��b)y�r�/ԛ)]l� `�-��p�~��4���W(�P=��B&���W��>q�9({
���joy���,%�3_>^�dV��;��8�'�K���gQA����єo�r��T��jU���k{G#�Z��C#5����͇u�eؖ�+��o�T��v)�_l@:�}ɣ���v�_xBe~��(-%����4�&&'W`���с}M�v�BGQ��UD���i�S�sLIjj��U����k�Z뿠W嫟䠁�k��OKO�Q����l�,�]e<F�n[{��0�}u7���W�#1}���yx=DBJ����<�d�&V�,������-p�g+�xvk�k�'��ƫ�:!�{� �+��;EОԄ�P�����^����~hqS�� � ���'�C�S�'�4�~hWsQ���j��#���#�����˾)F<���j:�u�*>r�8����7T���/36�T]kC�SW��{���AS^*��ή��Lp�� c�2��zJq�-mC�צý���s�jw~�������R�u��W2�(�%�l��--�qE[M��q	;c}�Q<��T����{À���v,Ș�ۖ�0mE65�h�"c.�n����%�|�v~8Y�w�^Iׄ��F?3bv��j��OPv��݋�͒�����P^۳gLw���4��qק�YY����[#T��������=���;:��JT�ɥ@��Iu-��D�]��7$mے[�t޲'Ӳ��oa�P���,��|��>�F|�� ��;{���<Ԫ��L��̂�4T�@�/0��ZJ�T�j��˚��Uq��f��2�=�D8d6�yx7��{ݨ-���W�:"��N�r1��INVH��*���%s���en^{U9�����u�����
�G��<ߚ,�M�R��S(�!�3�6��u�7�ߑ�Ui�='6J3K��Gko�?kXI�m1��	3����m�{%%i��nw��Q�Bx�QKj[+��4O1��N7��-��b���	)#/�^��#�%�r6�:64�rs���}�95k��/�Z�Ԥ��wf�dJ�\\�ƚ5��5T!1_95�=Bוeu( C�[a,��&�F���ɽX/g�Ҹ���*$��
e��rCbg K��+E���uڦ�����4`�]������jz�zU�vZ�YKY�c���U��o�z6�Z>� �v��+++L
�g����ɕ5�<^�
}$W48"�Jt�V�P�4�L��0��~�~�}�̪��Z�c6݊� �� ���͡��|ھ���Px��X�b��V�H�F!L����b��G����ngy��M�{{��O䀝�_jZ�^Y��6-=J�<�xfMXf��`��5�-苼�i�߿��H�/!+��H��V�6g�q����?���6�z��5w��WG�[Ͱƣ�M)�^�%�s�#1�	�ݦ�E��=h��U�m.( 箋)58ѕ�]ӽ�H���sd��=ճ�6s��Sd��{j�7��Oi�k�i��?����yR���qL	F�<
*2�	��0ٲ�'ڂ&{J�<�@ �X. I��@
��%|��^�v�RsOG=��s�@RTG.�����۳l_��nt_@D׷��a��=)%,d$�E,�SS����V;iƺ�M�|	K����e�����=n����j��!&�ݮ���A���ͷ�-u|_�I������R���Nj�C�ޥW�e��`8��8�HF[9z����i���[���@�<7��lj�f2�r��#�����`�+B梯��������:�ϊ�y���OB����:� �B�g�_��^�f�z�̓Lʦ�o1��ucc� �VC��.�*��r����𘏑�SR�t[m0��J���S��m����|:u�2��E���	�o�8oM:����t-T5�Xe�b��Q���Qt����~:��=}pS$�?�ꑾ�he�T~�&h�w����������?M��]7���֑'�si��Gp`K{��x�I�����BTW�Sp}�Ø讕��eJ`��zժE�L��GG��D�v��l�[�LY���8�V�����K.�[D)�l=�5�.�c���^�Α�s�����~��lj�z�`��E@L����g��oN˖�`�m�����[0����r��d�� ��D�f�Xe�
z�۵gU��G�!d��w=�����2\2��y�f0�&�/�̥�\�W���E��W�[h�1|@Ǵ��D��G��<�OH3S��?��̖4�VL��9T�@�ͮ|�E�}����}<����`�'�2�͒d�.e�=�m��"W��2
,f_cb�}�h�ε��G���n �	����q�I'��-������‭F�wL%��f�=�	`bC���^F�Tf��!�LO�,�j��puqQ���+���@����>�n1��'�O�\Q� �;��c�L����I�Q2�߸��6z�c�Ziǂ�
��|�kM���zkZ<Zt�od!�N��T�LKQY�Aw1����ӽ��	�
W���g�ڽ���V����h:�CtH�����P���W;�AS�ΐ�Ō7�]�pI���5$��YyLT[��rrR7D6�f��A�~>�do�i<��`C��5u���>�kA'��>:�4��*����m {���τ�N�X�<��a��9�S���S���[@�p��HyR�?�3�AO�U���}��k����2a��g�R�g�q>�z+�{I	�S��F���e��a;�ء!e�r����ꃒ3	-�ځ�gV��gc�2�Y!�j�[;��R�d�� �J�:�cT�S�Uz���G�����-�u!��	̋0'�Ѕ8�Ȟ���g���7��2A<�_�K�F�^������ކA�#<?+h�E�6�ج��ĸ��Q߬����l;H�f�t�T6"c%�ܰ�>�f��N�s�.5B.�m� Mi+4�u��@��`,�;����Ճ�e�g�G�o�'*J�ݑ�U�=�<��?��Z�	j�$��os����F-.A���J���/�;ܺ}$���t���A��6uL��pn�����i�b�w�C�]�o�E���: ��!Ic(K"��~Z^g�'J}��#o����""!Q���;]�ٳ~�֥���w�hٔ׭i��3|�0�[
���g��Myi��Bx����/M}�-����&%�s�F`Dm���M�l�k�٫�g���$w���犂�dl�Zū|���c����J�z�����W�I0ԗ�lW�̡¾sHRˡ�gD%{���ყ��KjZ��A}Mh�y�6�m�*��G݊��>�&[�x�.���V5ǆ���ӞgYƬ~n��þ����@��ЀQ#?)Q���W������?�C�*w��+>"��iT[��&r�$��q�k쵷���>XmR���-&s�����H��j���GBg!�S	+G*.ldK�P刏1��N���\k�Ā���<�AhI�|����QGW���gr�Jv�@a{��Mv���I!NLӫ �|�
q��W��^�ݭ�b����Fݥ5-h��_E݆AO�E)�S�q.OR��a�wC.H��L�0@�LF�h	����#ԹX���ܩ�7�7�+�kשZ�[��z����)���U��߯�@�euypnU�4F@r�c�:�q
	b���&V�$��_�j�-^�Z�P�k��}�ǆ�JU҂��y|��1�t̪Kau��dJLLT�v���Xh����s06t��z�u�|i�ALȾ������YC�u��?1���m�2y��*�<Wf��1![���>f��I)���Wnh�o���s����s��(3�'�0ClD{���0�Aj_�z1#�S�5��9��b�>=��{��v�-淉�}�ݻ�z�/�Y-����ӟ.�Rm���ә:'���;����'�5����>������m&�ʼ���0�̐����l�|
 ��Kr.�f��ؘ���﷧�,�!{��f�*,����k#�wA>d�;i?�S�o�������j�+�|�h.�S\1#\�Z�>:���[�}^�p�P�^�B�w96t\aqX���8��iKLC����΅�?紣�����{y(�seű�����󛣂�G1UmB��G�?���̚���=�')�EfW'Vm-�5�T`��
Y="�nii��k����b��\��5݉�*l{Qӄ����41���q��Ϡ6���[ob[�b[o��ZUz<s��_��樏a�,t�y{t��q��5��Qii�?�V��y�Fk��l�N����ni���f	C���1TA-}UK��7�h��8q��9����i���'xLD"�GަO�
�6oJ�k�L� Jz3$K>�]��%�E�V�l��8D[�9W�5y����-�u�u��+����p�����b�}����͝�R顂�ۦg�����K��K�T�\���7� ��g�p��1�#*����4�3�.��x�3�_�DD��򓭦��W��*n����#��M;_ƿ��U9t�f����9T-���>Xt�����E�sq�ݭڄ��7!&f8���bn(}�#���M1�g���L��O�t�ſ�]6�r�X������(��o��?v�X�n���/c?��.d�<E���Ƨw~�g:B}�������ܖ!kn�0d��,���0�.��@��esN��uF�����PͿ[���;W��%�/R-v��˽_�?<~����{$^��-����������6i��D�W����a�T�~�C��c��1���m���~5�6�_�o�͚� t�F��1bQi���y���>�N<:U��hxOǛΈ쵑H3�f�ٓ��gXGUa+o���)+�e�=D�_�ws~�(���ȇͭ^���!����M��>����Q!N������ �"�*����F�sl���y�Zvԯ��W1�nR�d�_)��6� �Mu��WyJ�Փ[]\K��I�Ei��f	Oa�L^}�3�y�l�Ĕ}I��Ѽ�E�ʬtx����?��;H����^~i��Z]���=�H5ʏZ�E|��(����T{�֑�[��!��
���VH�1�
7���� ڤ́��;^%��6�/f����|<�iuZ=^[XE��>V�ɍ�"݀��7��EwIb�1mO�����K h����:�5i��9^�E�:���߀�x4�m@�9����tL#H��f����~#�$�w��t�suph_�2گ1�I�c]��\L$ �5k�N�A�f 3"��sH�dpR�W�^h5�H�$�����������*�v;kv'`r:�����c��$abH�2-�x��x�"M�|>I�h_wÀ�G�q���E6��h5���v�����w/�������xRhp�$�����I���WVV���fw S;:;˥�����EZ2݂�"���RgL[忟.�Iz+�9�aL3��H�Њp�,�;��ɯw���O@��߆��9��NX��r��7zE>a�'K��b����:8+.abL*"$��k�^�E�W�/�<�&�zʀ��=֒!X/��c�'��rIgU�u��\���������$���Թ�Hl�Cs.:��D1h� `���x�PN���׆�����SQ��
�%��t��t1����7�z��v;廁��bL��R)�P�Mzdp؟�oS��EwG^�]��}���D.�C��R��G�=R�z�T#�)���iy{�L���1���Ec ���L���$�M�F�*XQ�%�Q���@W�Тq�jCx�t�I�"�P��\�$�?*���z2�#I��B]��E��t�%�t
����D~��h�8�Ӏ�E(��)�d�2�0UA��ܙR%W@/��хCC���0�C��dL�]��'Z��DF�R�(��-
���"�1�> е[@9���	�%E��N*�:�T��O���o�*����Ƀ��J�i��Ѫ?
Hv1�#<�C~Z�q��
�_��@
���r�G��NH��
��$�H&QXI'�|��l���M�!J��������@�j������V���_~��&7�\h��FO�#��Ph~+{�<FT(X���`�6��y�p K�s.�l��u�>��W}�\0����g�	�!y#�֍����z�u���@q�1r.�'G����K ><��T�U���#�!�-PT���n7g?!-�G�+z<�����m��[�L��G;�qsuN�8:��TW��\�,r�2c�"�F���5��˖�Ӑ��O�>n�r��%��t�K;�כ�:/��eh�<6/�^yIz���	��+�HY��¤@���΍K �.����R�A+C��4�+E^d\ɋ@�+��u����,Ћ|T�$e��;$6��S����j)#^u=�"���NE��O�`���+�nM�zT�I]<�)i+~}b��PK   ۍ�X��`H�  /  /   images/0b5b01e6-dad2-4c75-9695-e3d6481bcc1b.png�Wg4׷�!E1�P#bkQA�أT�W��(5BlbE�b�V�ZAK��ݪ�)��Zm��9�y>��}?�~�wν�������&j3��Г��1��h��e��x��k'����%:_k�������쯓�e�6�qA9�;�I�?�D9:�:K�������!#c&�j��|�}��P����w����&]��$a*
�t�*�\_�Ai��(�)KU#�C��[c5�� @�`BB�sh3oAA�È�f�O��d�.�>u�v�5;�?�?:ڨ�sn��ݔ�㢣g�~9�	� 4&������K����8`¨����8�)m���F�#������߰A6��槔)�>$��z��?i.�9rw=K��Li�N��qJ�@��`�Ai�)9�Ը+���lE+���R a�*c�	�����Y���?/�|��I�����i���L7��~X�Ӆ���_�R�j��[�� ��w��k&8
K3��i7
u����6�ܒ�J+�k7]iR'S3���Hh��yx�q&R��_�竱UVm����jq��<�ڀ�J$|af��Z���V���I����ݵ\�׌�@�r����_"�L��Y|3p�WUI��'�>�&�l���k�&�5��9X��@�;���y i����<�<ï�3��Mt�m�����Y=���G��{:n�3�\D�3��g�pB1����8���{�|g���&�h�+R�������y�+�	gJI��/M�D2���ɛs�?���WnGzܜ���V���
\0y�=t�q6���A�kh*��8ڥ���9cHlX�0�G�r�����M�pG�Џ�r9X@{X���~�����cY�_�j N0`;���L�~�*�8�&�1�W�)S�=�Si?T7�����e��I�v���*N9`��N~&E��Q�\�4�ɦ��ڠ�*m&#�b����:m��?(����`�]9��YDUf�Pun�7�N�t��Wqn��H����؜�W9��Y���>9̇�����g3������~**���JUKC%�5�^�g�\~RP�	+�!�r�ɬ˲����eL��-��P�I�|�K��Z��F�᫟�u���;�V�g���H�z�5�={����}{��S��PLjv��<2uڶ�@~-O�~8��uS�5�5�_L�Ycup#s��O�7w�s��w����SH���1�8�5,�GVF\��눱��G��5�<
_S������a��O�ӈ���BuC��^��[O3�O7%���F�� �����i����}��nD�p��<�Y��ͧ�vM��؈�4^�r�ӏ�E�)�v�K5y���|��ߧ�Y[K�P��q��g���o�Z �w~����;݆���bw+��?�{���{��K��t+����H`H�'h�z�;́ʰ>5���R�xA;>��+�C�2����iiM֦52�-��⬟+��X�[���b��r�5(��vc�?چ����.u��$��gos�"yj��8�Ӡ�qW��Y�I��H�&
ހ�\�1�[Z����N=(�@Qw�fvUO����K�:d�A�lv�wز��P��������;�~2�?�v;&�l/�q��xߠ"9]n�� b$�N:��؆=�I&�0b��pZK+<����$�\)4]@�Jl�
-N�;�év�Q{b�+.��(�20L!���#u�_�l{|v��

��]��˽�1��xֵ���
�9��YBu���$�n�wH�\o��LF�Cs1���!�^��j�JYE��`�z�x�r���<��BB�ڎ�J����}���)v�6Yտl$��kF�j4v�� ��^+�3	��pZ��Up/}�̽�����J��5
�X]���L�'+:/�w�܆�-Єw'r���"l������J��m�6?H�屺�����歶��w���|�����o��b������S,���/�uN�
�C�\kΗHc4z��`�` H=����.���&�jO����"rx��!J�<������3T���ɟX�Y���oK�?m�?��m_<�1�/����6o`;rh)�����(;`ӥ$��W��	S�T�<��]��v9��A?��Qd�`��f
����!/8�U83&�K �H.J��G�@����4m�D��G�"���hB>��Ԏ�>�%�J2y&�X�r����]�}�x��y}Z]�W��.�U6<ni�\�`&�v��Jl5K��i� ��Nj�}لF�9�k��d1�xi\Ͳ���j5�L�d'u����7�ԣ��.�T{#�5��MX'쬗3�Y4��u6H"DPS�h��R]���A��j�6vFd�f�*a�L䃥~v�S�{z�"��ur�Rzv���:"��MUE�W!b�d��G���5V���obM,����:�����c�uSfbL�V�,�#$����G�;ׯ	,:\zI��s�@d'&�++�*�]�o���[�`*��G]���$�|�A�:Z7� �����vrG*�<0��~T��鵽��@'QH�t"ĞW���u�U��9^�qg]����&���M�Wj�<4EtJ>x��"�L"p: �˷</�.�C��_�y�`���+��p�����Ou�(��p�Ȼ>��q�D;w?�j�i���쾾�#*�y�:�4A��7���(�lF���X+xn֘*+3���2`��np~��'>�]������ۺqi�iJ���c�F�<�ݐހ����w��zb�g�Uș��S��ŝ��N�P~�'�n�Q�'ْ����iG��P�8-�%���gwlG�+�v �e��fq�uF%�HA7>[ˎ�a��k[�u4l�g�
�(��I٪�҇Q�$Ј�c"W9��� w�4╇�ne7�*�q2^1�^�fE���^��@����b�")�䤃\Uw,6	̷�����2�f�ն���s�^����~��Yj�^z�fH5�7�A��Jٴ��}^}�ߪ�hW�7�w�u6%�my�t֝'.�����з�0f���ݩ���eÃ��9m��J��P��?�9�_H��'�S_����%�a<`��H��8f��Z�c%���0�f��s��J�f
��{ӝ�!@藵$<��l��=��zٿ��YC�[r_R�{�"�A,�;x~!Dn� @RZ�C��ɚ���Ɨ���"���K�Ѹ�P�MI#`�+���#���oa��>"��F����ػ�elGs�U���m,�����ۻ�/@��!�l���1��t3)B��j�%A^�V/w-�Y_��e�؀m�l�%��8�U�u?�	8/� ]wr��[\�0�D�R��а<��`�f�s�W�;��iF"�����	��@�A]�N�ߵ~6�e� ��J}������Ⲳ���	hh��@.l.ho�i�0b�wNE�K�>ǔ�_)>�*Ǳ6�M�eJ1^,����]��3����C�S�c^�â��\�e�Sg�jL�\�|M����j��"Z��ԎJ�BX�=��8��T=T��z�L��A�Q�T_��'�\����V-�� K-;q:�/��������C#+\���j���-VELv�Z��IkĄ���/Q]�Q�－��3DJB�J��Da\�A/����-�����1��4���3e�.	~?EYԡozK_'>N v?�$�x�ã�Sz_6��Q�;�0�zD�.��NQ�kn�ĳ���r��������&���},�ᅉ�lO��~~;�/@�6�C�" :ܑ젂���A�ޜ�|��z4����D���00Rj0�=���#@�-����O�>�d�Z��u��PK   ۍ�XK�`��  � /   images/1a17dab1-c3c5-4679-bc59-2ce04d496e8a.png��?���?�N��*ZEZ���ڪ��wP1Z���[�-���Z��DI���D)ZZj��� �� �}�����������yx��9�u=���:�55�9s��$  8���i  �G�g}cbN��q�_]ϒ�e��cX���}� }=�9��fi���b��M������G~.���`i7/�G>.��~��T~ �2@O�eH���/����q�<������%�\�C�O!����*����q����]�$�\��UH�^����F��C�_�^���>w�!�C��m�W���]�sg��P+k�o�p���Kf��r��X2n����N�_J�_4ٙR<�����k���oë����R�י;f�Wd�^��0_���B���ف�DL�?��H��1"�*����+�H.�/��E��0ڟ᤿���^���g������%*2�o�A����W~�e�c}�:�� k��og�  v[���
��ϥ~�f�l|�G���B� L�\��0�ARK�ej́�R��q�U��3�Λ�6�u�.��U�x����$p9�z�xG�$���º�� D�)�&��� WCc}&G;J$`h0d�h��޻�lO���u1����8��Jipp?!�#��͖�C.9Ƈ-]
�	F�Ó8���ϟz���0�ؠ5m	b�G���M��f%].f|腤����U��?g܆V�̜ȿ���q��R�T�3�>oͣ���|Na]� �o��0���u�S�n�HW�� �l�qUk����j��SJ�(�0*�a|c�ieuTrZ//H��H�D.��C��ϳ��Vg� ��+rW�QJ��#ԙ[��a;���f�y��vI0-ԏ�5X��?�Wd���g1�:���y�\;+�H}�sQ���ݷgU���c����� �������po ���?�&�m��dp�i;+�����9��:q�?Sy��L�m-�	,�F���=�KE6-��.�syW���e8]d��Ȟ�����`o���|��Yh��A:�&	��1��%�n:�5��W�B�n@�bF�u�v�	�\g������Ei1�0 ��wه��j�ml�rWT4�:-Z��;��k��~��BZ�ޕ%Uhn��8��5�C'f��5ӅW_h6�:��������3��@ȻW*t�+΀y:�F�ƒ�ٸX9�\l���@3���S;*�&ZOO�<M�Vq��>Tk®�R#ۼ9$�࣭^�$�Q���q�*��k?�� ��4R*����j>K`t����|���B�M1(m4�f�\I��	c 
�@<�u��N�x�\��ַ��1R+�}8���!N��H+ZW��ni芔�_�b)q��������!��c��ʔ_��
 (���4���u�OW{��<i�ْ�ƒR��kyO�x�"7iѢ��֠�=�46�Ms�Q��Iu�Vl9�h�M�z��!XN�ꃦ�8۠���8FK��Mb�+e;�G���,�1�?�������n��i"t �M�,0r��)�3
cN|�+Y�n�ڲE{�d�;v�����W�菠Vg��%j�[�T����?"V}v��G�N�U��ɗ?ˋLq*|�nv �-<������+�*'����G�,o��6ʽ�h;�=�����\���!�_ȡ��j��JvLK�J���Ш�*{��v��t�{��0��h������_��ed�=yͯ�Ǣi���fF�k�5~oSF�o�{� Yr��<D�m��v>��q�Ɔ��ٯ���O٢+���_r�'k�ߥ	�a�ޒ�vv3��@9�A�s���`�I���Qz<eR�dCk��A�$�,�L��1qx+/�
��SC;*I���v
��S�I�5�	�ݮ��6�+���Z����|�����\Q8�=����������ݴ�~#8L�:�Jߧ�)���Y�E� �BN�������d<�{?���o��H���\u�|[_%�ք�s���y��^��������E�8��Tkd¸�4��Z��ؑ��
�É3=u���ƥOa�)��-RȚ��' `�t�����=�,4�����N.���0��`w���hzD��CY�>6#��]K�qԭ[��'c~Z>��A�ƀ�_4B��Xpk>�DP7BR�۪�{�VQ�k{n�ޏߜ&�"<p�  r�
:��ϰ��]Z�Ju�k[�n�j2��.�E�ɽ��##'[8蚋f�:�E���ΘS	a��+ulT�N�H�tÈ��\a��3l6Y~�\>� hJ�mQP�*J��XAL�07��9�����ٰn����!�%�BzJ��?�x�*���l�?$�G�&��K9���.��p@���ks��&��+s_��r#���޹.�7���]"
ۢ�2����^m�/�v�k;U�=_��$�T>�8����FXX�E��R8A��஻=�b*��N�x�r���V#t��n�9���*`����S,�Y�z�-��-�����u�{I����0����� �����Յ).�/�$
����x����-�l�x��5M��:Zԇ�����ڈ"��5��GI*I�-�?�, ��bH0c�{��ڟ��\9���y�,𹲣CbB{²{�����27�C�zV�ue��h��sE��\�==�e��rb~�Vm�?˕+$����Z��I�����봑��$-e�<R��蕆��"��+���nd�a�]m#q#�]��N�9� ��N��vۈ�^I��S�y��S������TLo�aNQNy����\�kr`ɨ��+�A��s}���	z5:K������cD�\+��gs�V�3������#��U���l��X��	�UFIY�`^h[�����������!liQ�� Uػ����>-h�]{� �S =S]y+X��;�Wa�o�� �;䒼�2Kl�]���gVg�{VG�gQ8j� �.���oy�kI���+Z��k���4'�Q�d��R��\�q��ء��;�is��vs>����G|����->x~�]R1�rL�:��c�V�Á��'%�m��%���T�s|��*�謶v�3@�\)�� Ӆ��Ad�m�R�,��a�UTP��Ր>�Q�;�}&�V�J���]R	������C��ؔ�'mR��q���2�`���V..p�z�n�5vS��7�n�`/�]�fg}�w�Rv�xL��������	�)�E����ci���5��q�����`�����ۻ����^�Xc"� A�H�G�~3��J�<P!0jȎ��v��l(���`�}"s�Ҥ�����+ W ;��о�U���k<���1��~����cO���u|w����]� *����;�L�Q,.�s��Ѻ���W��K$_7��ު��Mi�l�&T�:�kp����l#w�/+�FmSȃ�/�9ܬ����츁)ލ�h?����L/Qla��3�l�;���/�fLa�/�Km'L��qS)��}����������O��
2 �;���]ϓ��q8���8zڪa\"/׸}�JZ�> ��	�/;��9�S����? ��PJS����s�LW�����m���8�b�1��HV���,= �����8[�!����f!�M'B��v
���(�$ӿbiI}���a��*h��&p��RX�d{��Bww�,7VB]��iB���t2�a��bV��Z�	'X	���j�Y^c�H(�향U�3t�~��:�F*)>ޜs��-Q�a�$�����m��T��z���o��Ϫ���[��X^
1��k����� �?�,��] Ɔ�m�������a>���)X�Q�l�=@U�G<�I�`����*Ī��)�G[�kޒ�r�U��xi
�!-*g�mEc�(㒷޶���J!Pg�Dj����+o�� 6KY�:��j�j�a�������(��Yv{�t�S�}�㜈YdU�Щx-xG>���-��_}x���M�c�XY�^S�m�T�~�kvaPm���w
�ub�Ić�cK��6)r�t�g�/ן0+LN��p({]8�=P��ħ��&ksg#��_���iWPn�f ^��w{7r/���s�U����n�V�ic���WMj�-v�eE���O��&��
��dj�,�{�y�+BJ�8��A��ܻ^!��"�)�J��7���c�{*-����8y�x�2��o�%3��:�uŇm���AK<n�����J`w~�#��@YT�Ǎ�%%_����1 ���(Ya�m���$4��	��� a��v��E0_��2��m�a�ߺe�v6~a��?�?W���.җ��N����g��@�6�dFm�6���(G՝��9����j�+����v&�����3+Z-����4*�:T�c�¥$�-�@��sK̽�͙����9h��4�:���;�Ƥ\#����y�Q%��j���X�i��5���x�g�5됥�h�С�ۻM�^��Κ�I�q�%Go�'T�
D�s���6o{~96�Z�*�l�9�v>��>2��&��ĩ�Q��7�f��!zDA���Y����|"%W��j�_��5��3�9nk�#�����޹�����[#��-��ȳr�1ZM����W��,�&�Xr����90rw�+��;�rɘ�N��ȁ�8ힸx��9A�ô�8+d�O��������Xa�#�kV��rT�&�z(�R$%>�
S�K���~m:^j��;XV�����ږ�%$!"R�@��x��%��=��Va>���8���&����^T���w�����3վ�����mw�(�V��nÈ�E����D�w�@J�A��������F~v'}��F���=gl݉��
dEBr��L|ɩ]ˬ�H!<Ӊ����Q�UL��_� {�_ͫ��h��-w�����<��G�c%#�x�2[+�"K�N��Н�KIk�N�EPe
~j��P��k`��bS9�Y6��&}���[�5�J~��/zp���1��oun�O�Z���Ѝ��a	Y�&�	J�����<��+ə~��5_��P�@_��Z���)�X��X��_��:�aJƀ��/X�lDEΣ��0ޏ��Sv䌶�K�S^��Xܸ�Tͦ��j���k~�U38��#.�hk��x�,*^EO~�S�4R����Wx�%���,6WUc7��_��BF����(�n)��&��\����Vu��&ot��j�B�]H0w�E#�4u��Xu��\.!��Wc��M�9�$�h9��(�{Ru�烞fԜW��+�L�ݦ���´|�L�-E}!��n�&�'�bn�(e�ǨI���� �t�	��L��X�LF���֗�J
��S^u9!:���������m�?�G��mO8?�5f��5|�op�QѪX�-Lg���	^�ٶ��6U)���NdC%��������&s^�P��S7�dt9�����&���ݒ.k�k_�]�2V6T��}
�ߧ��q�x+6���kK�!�&g��y����X�w��5��-���vB�.B�b��ry@��H���X8v8��q���y�g�����B���S�eJ/ǲ�E�I�+��;'㟴���2ب�T{�$�I�K�C�_���}r���3��Qb����}�̨���U���a�f����5�1D�|��|�z�u��ȅ�J�>��Pͮ
�4�=��������bQ��B=B�9��`9*.ZQb�ݭ��`{�>"��֮h�� �VU��N)-Q&��Q���;&uC A�`����_njo��V#;�0FE�&�oN׏I�J	�蒜֒hTU�ۏC('��qr��j��YĤG�UE�ɲ-7��jC֎B�"Abz���i�1	ŒS�R]�&RX(Mѯ�TlN��a�G!���p�o4�2�6I��0�.�x�G�-��N�h��EI���\�gmw&�ak�z�1� �4_XظjSr5:�Rn���[@_&����C6����g��l�o���?���V�7������H�'&�p�z�A�V�xT��h|�i+�`�rv��*-d!2���GHJɊ���;�wC�N7@H�( ���1�KhD�%��ѽ���e"���z��#��^���+�O�`�f`�,|�et`?�o��s�XA��j>	�bVs��`ě*hx����ݮ"��}� ����7���q�f���E�~�>�WY �޽v�Aym�̢�%���
4~�WA�3�N5.w~BkRE��,b4cM��ͫ�w¿�!�B�e�#q!8�/��Yb$y�M���~�)6j���4�XT��X��޼}��eP���Ctk���YA�Y��b@؅2�>�[��j��݄�0��i�a�Ǟ/��t<"�@�䖳ͣa�����埃MF�f}l����8��b�q�*�n�,b~$)�c)��%�%���;�/T6��	t�<�٧\4����GSw&�s�i�?(��_�l��H�ڤٷ��gVk"���7��:��nH��p�r��fd��&�7m|�s��*��[w��uB��V�����u���k[<���ʈӇ��4k}> Ws�c�>��'G�Ჸ��D��V������v,8�)�t�1SBdd�`K"E�����sMp$#�����AE3ݭQ)f?Eo�G���n3^��L7��㽐��*�(Y���P�{�_>ۥ�����u�/�W����l����>t]%��;�/ъғ����)߼6�����`�(�LK U���w'C�pF�DO�j��p4��mKT�ݝ}涶�d��d�_m[��3�����T���_�ʳy �� �f�9��ԙLn} 	�3�t��Fg	���z���_Jh��l���im�7��1����Z�g��b�_v�]�9�柄jSj�P���~��J����`��=�wd\TO��@Й��G��P�g�����e�d� 
��p�76���6��POFj1��"�۵pG�:x`�M�H}��>;����h��П+b�f���u�#ϓ*�{��|�y �"}�����B��~�������������ڜ��� 7����#�<�o���h*�5ȼI�'{^w�|D�KKČ*� rTOb�:���6��l��f�	F�P{#�"�8:1��a�){[��&��%YHsJ���:dx�У�X��#E����vA-0�k0�/�A�A�P�Èy29!���.�}_`*����Z7ѳ��G�`��R+����i?��,��}�o��l]i�n���S{$bǰF_ I��t����:E;h�_�ya�������R���7��u���:c�������{�L�:�AT�4��q&*�oh��l�!ۗ�e���oP��}_��7�g�4]Z��Q���K~��p���4n=˝�U�#�%'«z4�����׎̇�d���+�����e�)���Ӛ��D�e����c��C�V�֎ݣ�R�۩z+�?õ���Y�#�y�&��L��� i��[�e�Ͳ� �#��'�v���j��aw���+=�yC/���Ā�)�-(�z�
Tb�)*��/(��ې>�͠�X�
�:��/����/�:���
h+}Z61�M�b��@Y²�l���_����?��0��${	��O�f�7X���+��sm�N�;��+K��f�Æ��f�FE�ʵ3�܂�m�K�mZ���"��푷�L��T����G>��U��zV֔�.�~���V�ai��]�i+����Tv�i��r���s�rb�Q#M��>�0�x�j���ʗ�]*�̬�-Ǽ�eU��Q��{��cv���O����}Fk�~��j��z�?��k������(3w������eYΘ�ȋ{"�W�2� &nl��m��m�R��ă�aQ��U[��@�����+�W�kv�oMCS�b�sJؖ�B�S�=�n�t��U�#������>��~�4_�yA�%]�Z�~m;�^_mO<&�Y�~��&n?���ŅC������ĂzX�3�
��� �0Ƴ���Π���Q�=��}�@O�<d�,�(ƛ�Zݐ绔:���,�8�G�
A |���ν�YHԃ��=d��j��c�A*��~�5��D����b��,Hx���ul4/� ��
��-+��.�ua���v�/��/+Lp���������g���e�"eK\Ӓf��I^���[�̈��	��3\�.6C�A���vpq�3b�tb�J�q]q�7n�*�'<x�x�36z��L�����xPψ��U�ƧmO���t�����ݓ���.���K.&�|���3Y�&T�2�}��,�,xk|TM�G���Z%픋�
��o� {0��J��SQe�{��ц��Ɵ��2�=�൫(�H��4�Ki��7�׽̘M�7l荚�?xBcM���{r�N�G�nDy�jm�vP��]��!)"j�B�j�bČ��O�S��78�e�G_��rw��v�C��������ːW 	\"`J^�����"�:ƾ�N4sP��R=��YJ��=t�^�6+��G���i�{}U��bk�s��'�(%��ݖ2e���������wV�N��C}J«��q�����j�3ܦg���N����6a�_���	=�g����Fs@*5�k�	FÉ�v��{v�ch�(*�=y�c��hW�}��ſ��歪e�	��G���|��oK�/����[2�07��|�"7�ң���7��K�ȳ��r���U F|$tI(�t	�����xn-i�3����U�>1�\}����aF�7����U_������.+��ؚ��;ئn=����c�sNS��|��b�^��kw:V��V��m߫�b�3�৭��.��ǡ�P��v�2}�<�y�*^?��z��;��*����^��l>V��
���f�;�ʌ},L��f��_qྭ���4�-��8В�?ّm�F��2��G"8��9]4�5�o5Ǜ��Ɓ��G�e��s �S�����.R��4�cS��d ��.�6'$l
}����s�?�t>J��q����"�2_N�e©/�.n��mPְ%+w[�]Y�eCͿ8��Y��2obw��'���1b�O�2(����k��<��a���~Z���f����ϐʽ���C��W2�I�@5���e���J�:�*_�u����tF���OsJM)�Ih`�j��މ� ���\����bܭ��5����R2�C^���Z8GA���4��$��W��`�Ѹ*�"v�?�*��V�
�tL�Tଜfs힘G1������k��T���'H}6��z�i���8���������|_C$}�S����n�a�D��^�\�)�ԨZ�|�}�Hh����~��p�b���2&�te1f@�ǻ4�_hM�:���&��
a��&��F���JD�(�S�+���R�|���,���_�P��d���"l���lՔ�&�~8x����:�j���>�z�)Y�1K�c{̛\�{��s�2���X�4<�`�w%0g�N�?���N)eόF��4kNPj�-�,F{��B֩�ߑL����0eS�@�&�(�o]o����Q�r3���R`%?�x�P�a~}�Š��mh1�o1z�D[�8��,�'=�0�yQk}�	!%\��f��9t�፣u�(-9�ba?͌,���wka:����ŉ�MV�x]���4�:v��3z�� �-�}S�Q6�aܸ`)�$���#�p	ɟ疰%��$�I޾6
�砣�,�}�`��<��ɨī0���R�'k�z��w99.�&S8"�f�gz�9�:�$Z2�QL:�w���2��[sk�H��5�m��3e�D��D����~7���t'�
��W���]���wa%^�a����ϨHѸB �'��c7�YY����7"MJL���<�\�O�4��^�����w@������	��U�܆� �ث��|�~�b_��8�@�1��u���h��쒰�D�����6sU�����<�US�ϯ�>��&
Vqm�x�X�*T��j�ʳ��Z!r�H���ٺ#|��<����ʘ�Ϧ�ʠT�{^ό�\%���h��R�k��a�.�n�W7���^TGR�&��mѓ7"�[���} �N�3�*w߲��W��b���`I���8�<Gp����<�0<�C�B����8�].������v'�HTn5��\����g�5������ n|s�x�U��6�HG`����i��J���ૃ� ��~`�����"e;o��w���13���h��pY�3x�tm������L��hY>�/����+?�4a�C���������#b�2?�߷���`�<])w{�,�k�i��>=�7�G~G|XtQ�c<�D�e��������7ь����Ҁ��6�}/��.w�|��Ċ���J�	G�>�3R5R���S來,��^;�.W�8`���"ޏ\L$��?a{�N� |p�1ǤOC)2Pu�@7I�|����!�~���s���� yR;�����^+��.��)�)�ϵ:s8tN��T��и�B�ꅋ�G�>*�?
/E��/�U�gR�?le����\��؍*�����A�0�b{�����Iv���7s�IH�u�����D淄:�it~�8�![��+���f�yHc�=�~%�j#/Tn?i�/O`u9Y��Lղxq��A��*���t��a�"
ր%�1��y�K
?�LP��X��er�*� �|��
,�0�V�PL
x��Z�-����W+�w�Ǘ�d��'�ck6�(Y��-���<�]�^	�դY����)������
U~R�O���;�_�k�:WyB~&;�7.S�r��3b�����E����W`m� ���!P*q������u��Z�^���ӥ�c,<��?=E��l���P)T��[�o�������'wh�o%`����1��O�b?�!nJ�X��q���p�+�U0~g��kۑ���@\ߑ J�-���zh��g&&��t
dm�s����J�k3���!�j5I���>���?z�{#o��%�2�m�{��M�����<
�y����z����G����h˗�pۂ�=?�r���KrY���"�s_}h@�t��vB�^��k��百����yK��Bq�+C�f�)�8+�1�δq,-Kn�Բ,2�����;�OWNA�8�Y�l'�j��N�R,E��yv5"{�=��g��`An�Ȅ�ŀ� LY�5ew+�s �]���B1�y|�ym��:d@}Y�IB����i���7�)އ��������b^��؍�����	�}<��p�"p����-a۱��&���UB*�����)繦��V_�[����P����q	OU>�զ�Ȓ�N�xhJlB�Vk�����^W��ޒs~�ba��d)`Vpl/AV�15IߣX��)2�ۆ|�G���i���P�¼��S�D��H@�PX�=ZI�#�j��K�L���
��iV@la����=�cN0Fܟ6�Yid�X�XG>���p۝���s�`C���g�����Z�h�<�,���Vd����?�GU 6P,��.��j\t�OȠ�i!.��e�r­Xsm	4c(*�Z�sb�%�2�O�H������&+M�ed��o�A�%؍@[��Ţ�3�eg<������]ƪ��f�%v�{�Ǐ썗O+�F�;�F��:�ó�����,���$���j����徽�M��;iU�F���O��Y�^�(��n�0�;6M�r�XI��t�/>e�ҕ����q�*��QֽL��۷�JD�^=ۊ�S��~kk4����[b��0���'"�>BB�,X���ޘ���F)S����^^Y��e]I�N]y�",j�y�8�<C�:lN1;q[�I?��xϻ`����z�-�$��
�����b���l�2n�3�S{z�?DT�aw�U��p����ɣ�22PS�z��{�N��9��Ҥ�ᒱX���el4O��V��mV��T����e.����gfa!�(�4C+j�zzI���!Z���S� g���ݛ~�p�����N��ѝ«�P3���g����!�{��P���t��p ���Xg�D�pȝ@�ޞS�Z���fH��Z(�pEf3��w��O�`�;`~��������'��f�dG����i�<6TfN�3�|��}Ͽ�]�9J�]�	~������jDG�l�Fk��4�0%&RK���J�ǁ���z�h/�ޣ_���muB��lt����P?�5J�����6d_ ��jR�rd�{n����P��PO�����.�$����{���~	q�V�E����jp?5�q'b�,N��=O�ߟ>s�����s	/�����3��3�üF����Sl�E�>���	A߇�Jb>�3��J�� ����C��~�Q�����1"��:�%���P(G�令f�F��2����s����6mH��c7��<��(�e��B"e$0W�N|��H�s;���^�eS� R��T,�U$\����*��[����N��O�k��G"��I�!BN툁�C�=%�s�g򜹦		Z��Zx�k���1�����ߑ�Z{�i��T�����Oâ���B����T#_��;�S��=H�K��Z��*N^�k�>獠�/�:J��fd��[�	�Շ��U����B���?|�������#SR���:��y��Um��Ee�g��P1��EKt:z=�!�~�A��x�4����d:���/|��O�[�R:�H����s���
�����Fu=L�)��(��ra��jf�FֆDbǵ�6p��_�_�ὗ.TM�)�	vA���Dͪ���
�h�`��ߪg�7b�^��_n�0}�	���J�ڠx�0�L��W@��"��{�a��vvX,�� d>gKvQ��YD��Le�X`R7T�e�a�w��~	8x��Q�k�����o�In��Ϻv�"�-Rq��#J��''[���6�2��9�V�c��k)>�)�E&͊�_C'^�[�F����C��Q�p���j��̂����EU�`I�!��Řj��1A�]�3-�ck-&y!֘c`�iA��F(�+����e����l�H��Fփ~���Nq���ӱ7.+��
�d�������:�jN�ñ`f>�y
v�Ֆ�$@�i���d�,�����$�)8�r�(�c�G$�!�4���XT���OS������_���Z[!D��?42i�! s��ܱ;��C�\�g懏�Ju��F赵%��p^�9��OU4>���m�w��L���֑Vw38������j,�o�����@g��&���h�F��8��v_�f[�GW�|�|& ������L��/�/�z{��T�6�<?b��")�ޢu�m?�)�+b~)�n�w��n3_�?Su�$ܙ��-?h��U2�2%�wG�u�U��ax�s��ר%FA�m�i��-24h)��4��k{W꙯z�׊�4�d�`�tQ������ᡇ�܌^Խ�����SoQ��ڿpm'GH�♬i3,�2���p#�L�\�K����k,Z�T��4��p�b�7F<�lv����M��?3������9x2���O0z8����6�d�	%SL�r����J�~F�?Z�p�?��u���#+:��e��>��1X��>�rİ��<r�R��� 'a��Kj��==dB�O���d���M�/x��}Tl�ecJH��$�As�\ܒ� z�����f
�r<,��3� O��szk�oprg�uZ졳]*tPm��\��A�#�PA4��[x��G����_{}VE�'%Fx�|��C��x��s,� ���8���/� Z�D��Gҩ��}�*�̵�l[IU�1飫_��������j�E�,��Ⱥ*�:��su�W5Kjg�e�G}�&{V���/��)�(�܏��r��%�׊���SCŞz�e�<�����`��/�|�|�l����ƺ�Z�G*��|��l��p\���|.���]/�m/�Y9N�ն����/�������������;*���ˏ*��Mt^���(��CD��Ә�l�h�5:���ƚ亮��̝�:ȱ���Sy���߾���o�[+��e�x��ƸT
�9���_s(7��i�|�b�R+c/�C��O�ye>GŒw&����
R��?|�ar��l�M4YV�z]@l�-��q�&�u)rZlJ���9�fO���.���c$~���UQOC�l
`��wj�.��_ߨ�pɑT����I��S6za#��W�W
f��`�y�S2�g��֒��jii��?;b���O= �hSL�{�Z�+��x���!��ܯ����{����8��1���V�[�#��1\�T�ڴ��t���o�a�d�������+n��̷�;�~�i,L���y�S��	���y,�bwjM������Ɯ�+#��=Lۨ��R�w�8�;ng߳t��ޙk�Y~�d/p��a��v�e����� ��3�1�~�P�K����'����<>���u;B��6d�V�H:.�!S�]μ�(��^���A]�N����6KA���Ġ
�D+j�i��}�p���V�,��B.����~]��K���m��)�/Y@a��jmz�j2�	·9�vF� uN�&��͍Vu�]������� <�U�9ٚ���̨�/�W:]טs�(s2s4a��K|S�����;����?!a�9{�]z�⟌3U���k�l����0��S�W4�ݹ�E)g��<����Z�θC>�3y�m�K��N9jxRH�ۻ��<��ϳU���M]|��e��l�NZ˞����Gc�zu4g?�5{^{��8R#Ġ��&{��j�[��Ѷ���l�e�
Z���B��>�4�<�}�-�E)�o���7yЧ
�ɽDGc�<aj�<��"�S"����kt����k3�~����uܟ�;�� �U\i֛���3a�'2�ol3xc��X�i��[�7��Q�ĝsEcJ��Η|?r����Yʥ� �Y�P��u� ";���b`�/j�Y�l�|T�TO�uk�:S��c�7n�h�W�8L͕��l�M���B�4��O	�	���d���������|w�P�g��㏑�4,�1���Kv@��[d;N�ϙ�� A)*@V 3����)��.F�߭�0�`��S��8�Rެ���g���f���(�I�91T��p{���8
jK��Z��ߚ�PW�/�m�a������W�8�-��˩/��e��O7�s�V�� �V�On��mUf�t3��e�[���r��eI� @`�[��d�!uҙ�vQ�U�3���EJ�M)���2�{�ݑo�)���hRT��L\���������z=���;�Y3��k�B�����M1��1�#,�_snn���'���P�����:��O�˲�⿃�w�����A�������[h ]��h�.�|��8"S��"7�!0�o�򈁀&���v���Yv�V�˟?��fX�:�м<uy
P���t\�[�G����VV��Dc��e��t�ǔ��n���or�Xw}��y�����b�>���6�'P'�!��a�R��� �q�A$�$)��I%I�E�qǧV��3�0pHe�V��/b�?�ug���|�S)V��8*�Y|EضL}|Ȍ֊���'7N�!ܟ&�l��x����a|/�a���rε�77��|��Peh�Z�D��M����Dɶ��<��vEhE`Ӛ��<�p���0Ϲ���C�_V��N/-�u�)���c+���U��l�<Q��y	M��e̢0J�C����D֥m\x�J	�E;��b�eH��,�
��h]�X��c��}�e�����<���z�vwa����<��;�B��Fr��oH�K�1�����L�1���,(Wsn�Zd��G,�2� ��	JP\��2b�ټ�J�T���W��vxT²tE�%��~v���+ȞQ�w������Nr��	�|�f*�!B�J��[�� �ݳ����*��Q��S�Y��|���U.�}��8�#V�2�U�j���i�h��1ߠ���7nU�=g�^?+V��s#oڄ Ƌ�[5��;��7�He��Rd��&H��I��%C���;9��/y��S�w�FWO��,��{(��.Dw���u;C��i�_U)��+�Q��u�fL9��\W�8����9�FZzq(ٖ��}*���7�]�}��8ƵU��3�ݙs�&��f?P���%�B�ފ�����D�9�v��;�`��Zdk�G�'��%�_��!K��m�u��r�e���w
l��-����a����G>�D|��:[�ۑw��B�@Lib�ے.��oԷ��8h!O.�%NM8�N��:�쥖� Աo������NH >}�JU:��dsj�.�
��l��h�P�^�>��s�:��V���i�3��ޔo��z|[�|��n���Ďů%vGm�)5���cS�`׭N<R��<���L|�� �x��.��������$$���<���p��i<M�ƃ����Y���[��AH�#Q'��!��#ь���@�tgU�
}��!(f[���!L�^��	ʛ��j��H\ZD��h?L�DV�7qm��3#G�{(�\}1�4�z����;[���z(��2Fs&EUL��B*�ٓ��,G�Z�D��BkY˒���sg���RT�!EΡ9T��JR9�0BΧ9�I*��s69��ȱ��ad��y�~���w]�k���^��~ޏ���_ ��܌�(��N�G��#ߴ�:���?��gfQ1 �����p�"��	��)Py�]�"8/������@ƻ�o��5�����gy)&��A���y<#��ܚ&#�3C����;�Ȩ�,ݼD���4���H:���2�&
R0����ko� �ZF�W�����B��-���poш�^��݌#.�P�5[�zb�-�抂Y��n��y��?�oPZt�p[�����#��~AvXf�2�.K���w�+���%��F0�?����S��OU�𙈚9��\�֊����ǈ�HjG�7{�Z;=Q�FPi��!��"s,$�g�,�<\bx#���r��w+�������3*��p	���A���e��'�텸�N�B�4���/�h��^^B��|����r���-lH{8/?_6�rPc�p�Һ��l��V=�D[3��݃��l����S�g��>~��9��Mt]3*�y�2�NT0�R|n�bƧ��4�"#8���b���~���a�D�dZJ=I�o>����=
�k��)�G��>���=_�Q�қ�:�1���S���������!���#����0��A�qf�����ǣdo ���fGRG n/]�_�:��u���z�;����6S�
Tx=?��:d���u������k�i�ZB���dPi�:&|y��ܬQۤ}M]�����I�GLR7�{l����xv6[�2SN��]2*��=<	nԛaj�a��ԓ�cs��U�1�!�/k�@�RΦ�u-�h��-P^��-���P2'i��ܷ6��?��#9ɰe����cC�y��v�]N~��
|p�r,uq��
%~KK��2d�Ap�U�B��U"�f}�� V��*��?3#ŝ��~���aI����8��o~�}�@N�E��ݸˁ�<_I?Ϣ9���&���D�{q���w�<zITn�G5��f#DD]V�����BrF�|<	Nu�#�6��Lٛ:	�>	f�.�5��I�J��fOM�+Ն�(�~� �ƾ�-i*�o�d�F�� ]�䁫��Jb�n�'$��O&ݞ�R�]Ѧ:'R���[���-��%��	��L�kf~~�g����NG�u<\m
B�2x  �;�t�
����0��
��h����;���[6u}�[�q��S}���~����Jb����b��ҟV0�R�J{8c�p\�z6-����{������բa8y���`����T�I��cX���Qi�
��.L��G�b�f�oɶ{�1zQ��2����j�3�d<1k9e�}���G ��1S[֊��n�lDC8	ˠ:��s��L�7,��Z��\��ÑL� %����&'jn+��j0"�IjN�X�2{kHoT�f�?�|8H���.��n
�*j�V��*@w8��7����5h�D;Q|�y�������l:�a����9�+l��Gv"�N�ٞ�p}���*�ၵ#�k��r���%�*����IW}���5�<��6���E����@�S=d�H�U�n����]V�v�];+8*QR(��d����F����;�k������8�&x�f��x��"�l���f�Na�"Ͱz��[z�0�جA�����a�Ap'`k�E@uR�M)?t	���9��Jӂ�L_����T���w�QY�.1���O�ԌHOg�}6A�F蜱F�u�䣍x$aw!�+�f�[�-G�/}ZT-*@�*N��ݬԋO˺�t�4R��7f�n
KOv)�G���2�:y)zF?CW��0$��<��4�e�N02	��^����w��i�3M�m:e�MD�}Tŵ���8痤�IIj#���A ���8MщFb�g�k�r;&��q2\��ʦڇ�G� ��&��-@�d7=E�4|k�������r�m_��������Zl��⇚E5}����M�q��h�\l9���U]\��иweL���������@��Tܙ�j}U��!w�Ƌ�VK�����~Xx��-��B_�J����}��u�e���c���M���͒���pm4�j��_�I��|�4��bb�˒��b�e��̠�zݺ�	O�ي'.e�����Rq���f���.�d�4LuI\Wd�o��I���u��O�̖x|N����f���xy�3%�.~�J�������Ty]K��X��' 7:��h����T����8�͊o���E{����'��*��$6U{��_�P��Q!*�x��,EWo�T^k�k[â��VHns,۩� ����^��6-	
�8n�$s���y�d29
v$�W�yt�۝h'��<O׭�ȣ�'~���t��.l��#t���{��L������G纯��t.h#�J�T��{�%(wߧ^	ޗ�a�X��Bjt���,�n9l}X���D�s��S�*�R䛱�a�p�o�}R%�g]*�io�?�s�`*t���I��I��]9w!k�t�%KJ�d_dY�|ͯE#���u�;[���U���IF�@��&��ٔ|1�V7�[00�,����f�!X� m#�!椶 ��P���<�ٟ�DǼN�{VN��f���I�ʗ��Y��M�
�~��nC�`׀���USS���#��=�t��i�oND_AP������e�e����î�����7'�QN_,h3;���{t��P��N
T��|A��d����Ʋ�ۥ���ggb��@��<Y�N;@}r�@a���������/fj</�̀�]!�ٌ���Q�o��8���*ygi�����ً��S� �4#Au�7�p�\��f�g6x���Wկ���F|66/L��h�q�|�oy�pJ��Cr���$�n]͞�L�����5�A���{��:��X��R���H��	E�^�DO_�jM�_�O@ �Ծl��t�ȣ~q�"�,e����ƈ=x-�^��+_���5-�e���y?�}�{��pgr�R���Q0y�q+�U�n�\[��ory�:�;�<�_ͪ��k��[�L1���qk����5���	H�!J 0��^aIr	�-SZF=63püs��ق�mM	�G���M.4kp5�{��W�I.�����(yKz:#�(��z�(D�����sY�?�5�B����(���n	��Q��a+���k��⸲$��`��i��E��g�E�~����Ii��o���i�hCJo�	L���#�\/������v�e#>�]�?�H�]�JPY�\
T�J���1����pl3D=��Ț�q&&�=���9�,�.O\��-�\��9��o�b	��<%"c�u7 �������MEb�g.Kژ�~�� ?�������x6��?�RZ�~��a�;�J�3le� :�v�0$�
���R�`a���C&]a�<���G�pM�����S���z��>�l��5�Hm�G~X����o0Aq�N��U�A���}�G�iG��!)i1��$^Qp�/{T�gΆ��!�ʼ[��Џ�C��i\q-z������X��j�7͢��2!����q��L��
d{e��}zf&�@(uz9|{SI�N�Fah0�^�W��K�Nh�ܭ;KC<�x1��sb=�JVW�夨�_�U��ɷ������:1s��js�g���"lj��bR@@ך[ �{�v:	^�n�3 @���"��ݽRa�@	5�q�@�Us��x+L&��J���dN��6r_���`m'E�j�$�����Ϲ���ah���#h-ݱE�V�ӳ�{=���Q Ò��m��!ۢ��l%�˩��ku�������8�M7	���u�c�П�wb�y����pJ����Yݖ����~����M�5-�	�97x�} ��X_YA�		P�-��B���W2��|�������۩T���=X'`��-/j���C�<��I	�r-	��jP˳̧5T*[5�V���AE�Bv��c�6�^���/,I\�3>�3�mMl�J�y��
�YoU27��XS��G��ض�ŭ-1}g*�0�4���'_)׬�9LP���=7<O�9� 7��I;vmR�J#"��-9@�\�,̙^.u	�m�w���i��ڣi��7*�����tP���fkwz�lzV����.���y  ���u�\��K����@���T���:�Ѣ/&i|uO�����;�����t�F���Kz�ͺS�{�sQ{e�ӷj����h�����A�Z��۲Z��S�	��\�$��K��?s`�dP��'dW�r[U�Yդ�&3�����/K���{����˚>ϖ����L/ą��&�UN婄�6���������C4XI�w��ޫ�K�����SÝ0�"�8i}�6���/��΋�2RγY& ��	���ӧ���������7����"o���gi/�au�B�4�@��f(S�qCE��R��_ �\k� 
�"���|8��6���]Y�ĕb����qfK�jř��k� ��e����� �V1,a<Fie׼t&a��`�v5�Yip9��Q0��+����qf�iFP���D��ڲ�w�/�`��./��+���s8�HH�M�%&\k�U��c���s�\�6W��[�즾r�Jt�g�:�ut�n��Km��l7F�G�%��l^���.#&�� 6���+m��@�)���;-��/����̖���ȅf%xY�����2�i��6�3Y�n1����������&-MCӢ���F�b�ǣ.p����[���X.]�$U��S�-��ʾ|�mv�}���o��*5N����Xlz{�`�H��-\��t�r�<��^Dz
77��QX��TK���y�0�cd�uc�S�aU�Y�����S�)����A�&:=��w9�}(���'ⰚB�"|NQ	jW�M�~i�Ž����	�7�:��aO�W��z�Uv�*}�Vu�4_?u��DH��rh���`^'���?���d�fN����H�:�����}�z�����`G`��WV��eS<�~9r�ځ������38������+uя�; ���3�x?ێ8~o�z��UW6ԡR��=A��%�;]ϔ���ו�x��H��J�9����x}�l�َ#@��eGX֎{����$��P��s2ci���eNY����u"
Hy���v�8y��y�l�۷1?A%�ު:�:h��ں����hg6N���i�U	&������2����Y���	?XM��k}���xc�G�.��f^n��%^�%JF^Э��%�����vd�V��,T{�i����3�h����˱����\�q���~���]���z0�.�j��T��x�j"����}�F�� ��p����24j�{..��zڂ�~p��l�]R�kx����@Y���l�)lm$@I����}1vIQa<oiw���9�je�"�5>�{��} ���d�6�8Nǜ�L�I�{�N�����
�xy9.,����'Pݹ���h�Ze�HmA
q=���%(��aA�r��@h���걥Hp�
��H�U������`�����VR��h�Tr�����r�,g�NBfĞ�Q�`gsx�����o�vm:iU��3��}�JF�A!�"���zR�����;4���N݌:���g1?>J:�zA������a �
#�����;B�?�O��n��J��n�� ӷj;���t��Z��Rp4�vT�{�7���EF�:^�k$m^w���t�]���/&��5*�65	�Pn��Q������~3��V�0ea"Y����!�	c����V�>$�-�:�҃q���Z�Վ�~�ڡ{�cV�#1�Wدܣ�ͽ�Xn�����;�p���X���gC�<݉�F�эx^�%��p8Z���ƾ�PH��*��R� 2���EF0Kw����a`�o�DT��Y�}����#�#D�+N�G\�R�ᇢ���Gɭ6u�ʿTqݼ�����5���v����\�0����N�5�$���A8Ű��:7厞)�f��͸�N
Xzx� v`3|⚂ ���9����q@B���
����IL���/g���[ژh)��l�C����<9���e�7��V�>�P叭�[}�{�&;�|�W�հJ����&����g����g�K��Z�����as�t��>�����Q\��7D�����^m��O�n�Cf�"�����әL�n�S
e���xA�EKT}��R�ڍ��,X�tt�pc��w�z�~�Z��g��)�Ұ�T�z�&��2�X�w���b��%=���_J�������$�MՁ���/��x�
�SG�՟[�W�H�s[�kJ�)u���©�����w����ʪ����D�Ec �}H^����}w�修a�*
d[�n'&�/�$*!��˧��%����귯���TYB+��x�w�#��D�3+��Y����<
�U�dҺ*������U�׬qj�-������f���P%��2�Ey�ON�O�8��6��[�n�����D{�%&-�ɹ����3zkk/8�u��:�e��23��~�3��F�s�DA�#�jpe�{/D�}�L��9{3�I��LYG�S+錱Ƌ�.��.�,BχG?�/ǜsx��q^H��I-R��}��f�+�8+ͬXϒ/g^q����긲>�n[ڴF �
>Dn-iJ�sW.����9T�E<{��n��$,������ݲ�*�����B;���؞�Q8�ڣ���S�pCi綇�88�#6E�V�����z�j����;�bnI��3�5\��ƭ%�yލd	�K�[an������O.�ӹ+|��H����ϱP?��K?�(�ń���V�tDB�^CD���,�#r��S��]2��5Ҳ�� ?k2~�ҧ}rn�XP,���ݲ�Tg�j�O��
��G�/`"a擽�=���|�����-��G!�tr�mB�-��뷸���ش�g4�����Q�(y�/,6Lܖ�G#|��9O�䤤��u\@�!��ާ^APo��g�rqqEvjR�57�mF�ߒ�s�1��.|��?��4�ݡS��1>`��XR�eqz��.�2�I�ԯ��ڧ?=�u/s��<�C�=��/3��!��K�Rŝ�xQ��·����𱱚�,%��N�7�E�t �2H���ףq�N'��$R$���O+�r⌁|&`��|u�v�nc�D1Ѹ���$��p)��������32C�������8��a�-����Hwߛ��c����R��ʵ����<�F�Ɵ��Yl{�G��ɺ�4��x5��f����n�F�c������o�X�!��̼U�c��/����|5��i�x�������]��ֻ�2�b��7&����?��5�o�������d��}�)�(K�KP����<��U����5�+lhj�8���G#і#�Y�F�����p�!������i%�#���I0Kgk����b4�N��p�n�YZ�!F0D�~��=w����������]��^o=��.���.�88�(cc��x���x��h��#��:���Ѓͤ#m=%q����ݘ�<g��1�9��,�w+�a������V����bc�@D�?�΂�0Fɛ��K{��Q�3���.Z `�Rhy]��յ�}�TT�g`���b��5v*�^��}؜9�#�I}�|nkN����s��X�@!���xm? ê���{U(>U���
�+��n8MB�[Z݂�����,�}�{�A�E���Ȧ�S�3Q�w��_Y�����$w���|�&�s�A����)���KF�aK���֙�;���v��ϖ�ʋ�5j��VjF?'�!�.(��-@!xI��6\��G��[��Y��xx���!9�w����t=kp�*��iT��W����k\��7���b��22���F!eU��6&T@�&n�.��� ��g��ME�G�w�o8F�'t��5,>�Pb��L�n�����m�;	�9��3�c��±�y�N������Du]D�5���c�m\ub���G����Kvt�k�[.>Z^^n:���:��:n��)�"������>�\ʞ���vv]f�{������~�z�5�,��F�wn.���֑ۻ�Ϋ�j�I�F)���0���k�
�>�3��P�����<cR��-Nʶ-�nB�w��y�Z������l�d�k��X�J�9��ٺ0�-�*��7��*�m�z}�n�.�:^�U>����䏹��W��{[���^�R��8��t��^��FAw��"�b���Þ�~��q��m��C!�խ��|��`��0��X��3��`�1d��pA�]d���Zg�������U�{��9�M|�|w7|�*��^�8A�	�-���,�p�����\�U܇��~���4MFāI�M����l��#�I�:�!a�r6;{�����Cb�G0�F�|�4'ԏ2E#t��ci=	%�V�?��H��g���t��҉	�!�_�[���:���U(e�!�4d���!!��r��f�G1^VV�X�zyaF+c���|��"�i�()�zh�3l�QT�CÅ���!O���
vk�zn��1�42l��E�G7+>�t_i�8A�8Ş�0��Rw��e��` +��(�~�����pG���N�����hƋU�Q�O��_UGkΌ���(��7n���,�`d�>Śf~�\:��ONQ[�K$�W7;�ѷ&Y厊��7f��Rv��|Ir�p1zU͚is�&�o��T�+�(��=K;����%����Q��ȣ���T
�<N�OϷ;c$�C�w��"���-!+�o��V�A�i��owK���w`"2uH�E��9]�OQtB���08��^����o��hb|�#����mC�ѳf;Gk'uM�k�	n�$!�����{0�Z��1h	�u�l�(j��rù��,ڲ/'&/<5��Ϝ���)0Q�SW���<9���}�F�5r��e?�pz��IZ`�Qg紬E���/gE������9��`���F�)E�u�ae�{Nѵn:b���Z�r�)�MSCgn�x����"}7!�.=�?��3]�n#���C�l�Ex��֯ 9���������LÊ��+����=�˫SZTQ��[�z�v�:@\��co�rn���G�����\�Ղ�¥p��t�M�8�� Uq�j�����D�Yƀ��t��;�ъ��kw4�e�����'�F6�񴊊�9�ə�Ǟ[����_(�؍h�(�U�"[���÷F�@.C�ܷ@Y�C����c"�PDE3x��'���~܄X?Xrq2��[� ��Oa�J[on�pbo��-p��d�޿!�g�2�㤁�J�f�[ө�{��8�L���Ϗm�\���ڪ`��?�m�T�Y�ա���%��d WJ�3t���kꣅl��2��E�פ(d�@Z����F;Y���t,iy��Q�ad��*drG�u���Ak�u���K��A�������0��Mؤ���e��s��e�#�v���
|�vè�I��c��
.��Ft����O�Н��č�:_\V�,פ\�`� �_�����A<=��JW�H�T���'<܊k��p�B'}�B_�¬�?H<K���<����c��ް�w�Y�}�D:c���ș:��
.=��gtF�?�.� ���PF$�/wl_��i`�z�]�$�Ֆpi��]�e�R}}��ڽz���qr��I�%%E���^�^6��	�
��B@�K�~j֩��D&)ڣ#f�,�47�#w�-�����YqUn�����[)�W C]��%yr�]U�xs�A�$uҔ�Og;��K�L���*�x��&�]��p.�W?Ze'�x�\r!��B�P�B[�Ct�yS�W�t�����B���	�ˑ�	���q>ˮy$@
J�M�;��r���kl��TZ'�t�z��d���t�`=�v�AS�0��_{��u����p�ڙ� )й��&t�ҽ�/k�rk�ZM@�����(���v:�A�eg���X6Z�l��ħ4�v�u�G�G��d�r�������W
��|i�hjk9r��sXT�^L��xп��C�t��|��wH�Yۢ��n��j{���=P\�K�~�zh~�A�^cp�݄y�G����w�$V̦��V b�q>�Lĳ�J|����� )ˬ��IH����5����GC���\���
��Y���Mq-��GI �f#���Ԓ`,�gB�=�>���^���N|��_�zW�H!���0�-F������ڼ���ᓩ�sZ{��cc;腬�#��9�HS�Co��w���"c'z�Ѝ����N�9~E�A�
�0�O�P�TY�i;��sEi�]/GU��@_��	�B������G�������RE��]g��W�ab��JBt�^'�Û��(�<J��,p#��Fx��Jf��+�0*��7��f��{@�-�=���I��e��<��ڋ@����8�p��F�<vp1���t�K_%����ڤes�A '�(�Kԧa7Gf>���ˑ~��$�Blɒ����A�j>���x��ղ^�!�K-Ԧ���n�cO��,����Z*�EN��uSFFS.2���Q�I���;Wh���_���"�+<_ %�%�<�-���]���,�\*h���γۺ���z�}	�&��sP�J�c"��L��թ՜�Z��݅��~�\�k�Vv����4ͦy�齫�7vf�	���y���b�Ӣ�x�&8��{��EӖ��{����U�L���%AZ�A��ƚ�F&77�v��3�s���!�[������W��WvN�.y��XZ� �K�A��f����a�B�~�����)��a{�ݨ���P���_9M�8�(�ڗ�b�
�oֿ�:\M��� �%x�����e@��6�z��Ղ�� �-5��� u�>��\�M��y���LLS[�-�,�,rX�ΛC�M��:������ޯ�gz��OŦ�T4�؂���X�׈�閹?4mW�繽	��j��|��Nx�o�RmBk�`|b���:������yY[����Qrr�3l�.�nTA�s���Hz�	QQ3�����>�5ޞ�<H�oA�aܨ�m��e�%K��V*�u���ٌ��6Q܀�4����B,>=���(@K,G�u����\_K�[�W���}\��4�z_�HSEu�<VM��m��t�B�[E՝��U��66���Ҷ3\�U+f#�&��|�Ý� ��e�
�>P���	`��p��?c�]�m�����}��7��+�Z^8��U������ڼ�/��P�io�������C��+����u�����|TB˖�rY��#�oʠ��)�й�۷Eʻ�"eś;�"��څ����"ϱ���	���`�F�3��>�W?Y����}-K&IU��|U�%%t@;=HfTM�#�B�:Y��y���B�ɏ
� N3�����Q
��'��8���hG�lZ��(j䟚�OK�P��u���,���bCJ��˭�����B��i6,A�TϏN#���8����Bkۮf�'kb��7�?�*ͦ�� &��dH��5vH��}�{�9�*uj"�fk�$L��W}:���^�KA����{�Q�S�6y�H��*cT�SY6�sK�2eZ�,�'��ؓ.��wg������ur�0�LڌML���n��g�D�����=�H�=��CHg�dI�R��i�K��A3��`��6�����I/W������j�%���iFo�8�i�/����e�1ʪ��]�H[ԭA͸�9-ݕ;�
�>���Ŵ�HK�*����l��� �"��w�����`��֏�8�bmi� 5�lc�t���}����*�u��ay-���G]��J�of����"����F�0��z��c�W��F��I���U�m �5�D���%�i���;W9�}*�����'���JD���2i/oo�2p�!񓧯�f�e���;J�.���#i%�xMhX$$8�2��JJJ�:��&�*8�pǫn�N��A���Y���;i	��ҽ^a�ԉq\�]S}0Nj�y���ͦ%j)T���hd��%��Ҧ��ҶK� �_xLΛ]j^9��Yw�8��l�Р��`�[��Q�;Ot�����dY{��lU' xҺ�����W+x1\����$ho��)�bj�;�:qև\��]�7l욠|�#�W�\��4��]N�I��n&�|�Jg֗�p8�5��Q�7�$|���)��!�Uu�3O��ť1��l:�9Q�L��{�k:#-�l؃o3��b*�\�3�[�S�*���}���Ɨ�����h�}�C>�0پ:<��5r�7q񶓗o��)D��m�_���刜�e6�� e�Z�W��:!��אffî~��}�E^k]���6X��N�-��+�L�n��:���t#7WlZw��k��|=�#*��	����E�ב�������x��������r����̕���r�Mc��DN���^3n��ٕ��GTQANh�#5�\��7"���dp���F�
+Ҋ����֟,���-�X�:�'f;�DÕ�������~�����zU���.9hە��6Deimς'%�Oʥ�
m{�_y#�t��Ft�x�W��+'����úu+�Vu}�$�:��3p�WwJ>H*�>��3�I��G�Z�%�T#!N���Z�C���-������ӛ𜷰s?��)?��� �A���f���������Y��tNLH�˧�l��+uu.\24z��Xs���n�wr�۫��Ͷ�=���П5Mo�ۢ>u��-ʈ�����[?���ð�QY�#������8l�|)�f�
�&�H�q�d���1H3[��	]�$4a0[PL^
����\l��4�<�m�F��I���
ȷ���լ�i�1��r����4���\��%�9�aM�"-�� �w�+)\�\���{?^W~'�ʉ������DC�L���D����D{E��m
�;� �!<���=1������
 0����de�L������F���6�k�ט�Jb(�%3�7�k�EB�+*)E�o>V\R ���������0e�&��19�N��>[]��y�$-���Y��Uw�� �3F����1�7��U�m�'���4'�Y ��(�
��$��4��
��I�RM�&�ʻNoM���4�
-��m��ib/bǚ���R���	ӭ&4;��-|9-b*�y� ����S�V��Ht�U��_ψ�m�A�ޘY���g�Ag���6�.aw���uwӼ����@M�)-x����j}TA��@��9�}I�Λ�|�~���=���zT.KtEEŋ���ǲ�̑�/�q�&�g�B������C'���]��~w4</�B���*{�˷_nr^�m��1��PBX
*�>T\�P��k�KQYֲ�~Ql�����������n(�`�UM��	����,F܈仅60�̧&�־���.��bjjJK�*�Bcؖ�[�t��*�2u����'�l�L}�[	]��n�gB(�Zi�����L��;�B#�\���si��{/i>���\5�4]�Ȝ�|����� =�#�j�Xī$C�(ȵ,涄
4|� �?4x��j��}���ը�r,0���;���o���p���j�zg*�ky�!�m��I�4�~���.9w
�1]-�ܵ0Y"]�ؗ?\}���4z�]� �	�+�]j`| ���m�����1R�W�)`�LI��ƪo��8��ݪ}��A �ת�5UBAtE,<q��K�����Dl�FVb�l��@���\� ��:1��Dd-V��R�\3���8 �o���1�ٸ�cHO���rs�_���l�Uw�3Zl�O73��"���Z�q��x��eM�R|�+�ސ�-[8���(�~.Ϡ�y�J���g�U1÷Uk{��l����Coa:g�\8�v:r�C�;?0WQW#8�$]��7JN�?rA#��#��A`6��`�����l �]&\�{K8��|FM�n.��J��8Jq"���ȷ�飽V�r;���x}�r�=xJB0���+��{�1�ϴ�g~(�3�{U[O����ׯ�9Xқ��o6�oS�O|��R[ܽ�=,y/?�C?	+h\��O�Z`+sKޯ!nHƧ��"�A�����ǧ�#u�B=I��s7$�ߊ�D�=ݏ���,�/����I$�1�.����C. �L]��7�c������Y �00$����؀mU��/���Z3Ƌ�t�eA�3R�%ta˘��� �dh>V���y\�> ��qn��EiX��}Y��#�]�������A'8.�\���Z�t�,ܻ�cD2���Яb��̄\8��b//�Oc2�:����e���2ͺ[�io��]��¶���H�� V�O�����X���V��Q�2��/���F��W���]��	�,�cξ*�����$o-�3a�Pg`$/ˡJ�R�R�m�����Z>V%cs����P*����gwgssx�֭�Z��Z�p�qDp�A$uI�y�ݢ��<�>�O�7�����4�����u͘|�y>�fR�7����gLf�܉�:9�7���6�3�k6�����_��Ƈ?1���6Or=
���e1ߨг�v�T��vRl����j�N;������$�Y��B�D�.�Gk~o��c�mСn�:?%w�����"t�@݉����r��,~6@6�t|�q䮽�fc}�� 8b|T'۸���7��Ϳ(plQ7���+킂]�HߑY�e���`X՛|�����2K3����xß��nl3��Z|�W7%�(OS<�D����
:-�I�k��F�4%��BL���/H�9�7�:���qn�u�7\����v���{{��un�(g�?�Ť�.�$2n��~�1�+�
��7��݅�8�8h��n�����1{� L�g�g9:4�[6���*^
�f�q�,z[�����L��ԉ���e����e60������̴�HGz�4tY;:��0Gc`��0�M�ᠵ[�C�|I��1OފO����D*�|X��@�`|i����¬T��J�Q�r�~�n�n�'Ln�B�B�e�6�ZC�^
�<�8����OW^a��'�UW�<~hݚ���Z��������r��8�G8���G�L�"H��ʉ"����Ͱ�MU���|�W8��0��绥��'�У ������rW.ȁ���(N�\�@SLҜM�&d��\Q�V�l�԰���=_8z%��h��|v)< 2�s�����PH)O#k��仇$�Ћ�:9���~7'_Z"$�}�;6k3��d)H�J:�أF=lo/��!0OHo���Ĕ�}������_V���bc<�0P�("=�&y�u�6����=+�\�>KU��_.�VR�-���2��=�iӍ����-\�K���픬���~A盧�7M�9��́M #���>�VLZ���S*�mk�rX)�V��5�0��J���fΙ���ߑv���nAMm��x���U-���y��w^rG��y���h�ᙡ�ԟ�kU��2U�Շ�3Z���2�5j�p�ϖ���Hc�-D�7����L��05�'���!�u�w��Ⲓn�wBpR1�R|�rl�g�p��Kyxq��󐱊N��jA�����u�k��R��R����D�����^��c��̦*x�c-,t�x�Ƈ��ww�?��d�^�-�*s�mM�$�y�y�Q��a����G$ܥ+�C���p;='é�n��8i���b_םb��D�s2p��6�Gh0�裕(��L$�!:(`-M�dM�f�i��;��5�*���{ ٣�s0W�p��y8ޞ�)?6@\����|�oNW��X��!�D�	F��� VʟIF�E���&��Y\3h݄_#�Tll,��j�P����NzV?�d*� `�T�ڔ�ECc�9_f�LoL��7�B/��u_�O6"�̲x79x�.a9�Su���,���:k�=@�
����޳�|�T��jOK	[�<���=s�ͣ!sH��5���h��0Ie���VP�1�/��X
��jV��L�}|}#���営V��-sf�0+X�3VY0�k5���S8��$�B�Zl
����]����k�X^&.�W�a�ͩ��y��4k���O0ۮ�/�����s�� L���������K�u��1ɘ����wmt �FnN�R���7B��2i���Ho�F3	Ӽ@J!�I�����?������%������G������zs�`�J���Ϸَ��ol�����O�]I���$�Z[��S������:�T�Ьz�p����c���=��l�d�e�R9U>}˫�z>[
�&����[ۧfj�뚸Q�a�ˑ%YY껽Xw��#�A�:�����/�y_�F`���8��%�ȽWM�J��ɡ`����d=�3+|�hB'h��9�
[�����~�a�䳈�M���;%����^몯i��?�KOd�l
����A���s�+�%p1�Z�Z@*��'��p�������QMe��p�q,0ذPf@EA@�:� RF�� ��	 @,� -�4*"Ҥ� �H�D�HB�&�$����������w�����d]9��}�~�����ܫ�m�RG�%!V��qn������7YՃ�ǩ�y��0�0��nG��S�Ӌ.���|[��SZ����@��LX�u8>�u�x�o���{�v�~�@�`��MҦ��9N_Ī�m�K�d���a���hqx�5�b�;��3�����s���ۼ�E�XJ�H_�WOLV���'�+7Z�y��ܔ\^����Ϸ��4++��*�I+E"{�ƹQ�66O����?��-�F-)4�KT�r���Ӎ�8���ٞYjc�<r�����t�I�%�Ȩ!69�iT�����3���1E���r_����!��[�
/>�����ʮ荼�v��ΜC`����j����߈Cby/��g{X�7�Lj����T���[���z�*�'z
By�p��Nnni�Y��[�Y�^����J�3�W�-#�ȓDOy\�W�ZV��<TZZ0����255L&��7��OT��9�9�.����عleZW�9�R����Y��y�g����?�G���hk�^3riu]ގw�x�w�D$�`�������v�W�����Y������LM�y�Ҕjz+����K�����adה<k	ȣ^Nꭑ���z �?��ǧ�ɔ�Z����C��i,�0��&C�DO��������E}\X%�<F�3Q4F.^8��Yw5G�{���G���P�c�]����oj��ml�0IG̞h��r�l
Oߪ
���K�����,iU0�7���k�Y����>�A.��:۹�
����Ε�r�P�R۱�M�xuT��^���ck6��#Nj�,��F�����%{���z�@��E//DF*W?g�`"��%%��	�`UqBN�Vv�Ve?�+��lٞ���**zoV�.?���7���W�Ⴅ	�d��uo?��-;�NoM��|�R��j;?.��k��}�1��e���-0��n<9��t��Z}e=gYA��(��p�yJS�gi�#���2iG�Ȅ�g���M�]9˳�xX��Һpk��*}�2b� [rI�QZ�G��"ʍ>��mқbմ��|e=J�$�rN^c���<���Zs��P;fmh��O�)��vp7]k#���:�D/�I��?j�?�v��6�������9�8��1�7�����?�w�c��ޗ�3}f��L����
������f΁��;�\��pB.���ڗ!Y疪q�z>*�@�����#�/��)��	�[3�c\uA�k�u�]�A�X���:�Q�e��)Nd�E�U���z8�mfƝ�5����)���P��wʱ,o���4��E=YY����`
ɛ�L�K?H������s*�ď�����r�emJ�"�CY�X�ٓ'O�g�⡃aI�[�?G�n����a��r�_��hw��q�
!L}J7�H|������=�x��Ď=�l�(�K�/�U�A�$�1����[�����T��Dްט!Q1tvy� �gh�#1ۄn׸��C���F�.���m�n,�Mo��N�c�ry��b��� c�����K2�*��*���6���H&�M���t��m�C3��qx�X�� �аXF��N��#�[x��h�E��@��>��w��;��c0M�9��J�$�/l�e���{Q�jV���k�;{v����}�6��l�0�P6�X���]��@�}55Z-�Z��-=;���+CM�·?���̊v�z*�8�H>��_�D9�Ŭn�F��t9�)�8��V� �Rt�h�5٧�Q���Sub�c�����P�F�x��{�>�9���vmC��ͣ�y�� ud��/���I:���O׻�l����l�RY�_٦��|������?<�r�mL�rs%>�=����v�%������S���x��
����Of.���� �E���΋�
�	%eN���ote�w�,�ͩ�s�<���] ���|9'
Td�B��@��֞P^���n�@�Yz�@�B!���|�<+�L@�34����7J"���o�;wJ0�ӋUP�cp��!�z���X=^ʊ���w,��}쪠�܏�H�9��\5��o4�1N`eY������/_���@�P����csɑ}���7n�E��&�Ȯ7�&YQ�?�%ǝ{5�4L.�d���R�>�p6��7�.k�Q���Kkf��!>���L*�I
H~�Uٹ�iڵ��HK�d����a�&��}������Rs@l-��mI* )���`����$Mv�����<� R�=#{���t
�e�gO��S���Vt���P�:B��^��:�/��X���ʼ钨�����Կ˗�f8�%�5�?m�8!�t1F��Ű��H_;xϯa��@��o<��wPk�+Y���ݦ�D�O I'6T�ѧ:8�����g����?������p��][��u�O 
�Sۭ�$�3�?4Qy�Vk���m=h��M�j��U��{�(�!��fח��H����s��Ml~F�FG�tVɷ�ܗ��y��Q�A���(�����zb���z�)��w�T\������劎64QY��4	e�M!�/Bq�%W�_ױ�/���p<�*��P�7"=�CϜ��wFn�T�,EFl�J��~�&��x���k��nH� ����|�ʩ�����s������,ӗ#%SZ
��Q�v�Ȇ?8�]/�v<�_.�t:P���_��Y'�oZx={���\���x���!8zx�X1	��Z��4�f��uuG/խ��P�D�їf���&�j�L��y"3.�Ӣk����6%�͟iet�m��1�ȲϘ!�DeTO�c�|��_Nb�.�7���WaLKJ�N9�wNњN�{� ����(�u��yÇ*KZp�z>���G�:)��D&�oJ�@2T��zzͲpN1��"|���;�g�䱝KO�)�e��x��mu�B���3���(X���W�y\a�ˣO���I,q7OO�`�4'��[0�sŞ�Ɏ��^ﵡ�;<�?+����P�c��#�if���p�)�w�$�}U�;�LjQ#j��0�_���'������*��%��{��g��GcMU��z�5֩�W�~�$�SP��������ZC9���ew�� ���1�N=g�0���<NW����;P�ɹ���u��!���FHܹ�� ?9�Y��D+�{���qa�hI�E��qs�׆�Q�y#����ٕ�Q�5W��-G)�#-o�1�A��/�~�4P��a�{؋���ɜ�&|Ti���eQh�!��	GC��ɞ��2tDcE��LQg�B~�}g���c���ޒ�l��ł,5��԰���b�&�U��V45�`Nſo���}R�W=�����L%j0�GZ"��Uѻ����[~ik�o�hi]�b�ޟ٬��ᆅq��B�^��4y���uiQ��47�ގ���LY$gS?K��؛i��I��ȵ���I�0����O�MC_�߂'6d'�!�,�3�jSɘ%��֊o��F�ₕ�i��QQY#k
��������Nm�:ݱm�1a�V���{�t*k�v�2m��&h��O�0c�M�$�V�)a�3�7�� ���]���u]-l��N�*��Xy*��3�0�s$W�>�}�zg �p��'��~w��龠.Ul�;��Ҹ������Ǉ��U�*��S���	��r�rﴫ�^�)`�z9��5_�w���u|�v�~n��R6ݑ�X��-�iE���!��DFQdUg͒����U�o��@�	��w�Ʀ�X;@�_fff>�'G2�h�
����^+�).:��9�	~���3G%La]�6Q������������$*�t�dԈ&����i���9H�.~`O"ygF�Mb�F��-+����**àl��L�?�aXFE]A��$J/p�@Ԏ�$N�߄ƅ�2t4W)�M�#������MI�l�#�aR�x���0Xa�3n���B�T#s�^N�L���}V�t�@��WM�?H&=�9M�fIXi�#|?PG5M	�G޽���=*�7B-.B�A	�j��[�=����MA��{y�����jח
J`�g�V
y�L�P�5S6urvPgz��=Y=ro8�t��~[���%=���W���Q�\��U�ya��e6^&�ŉ��V�QV>��昧	n�pE��(�-��bȳjsl��G���b�J�.7��`>���Ko�&�&���z�E���C��O����r �����7��A2���Rl�g���G1�xpA*���3�V&^�\��z�o�6Ф��I�\�x�AKn$�`u�(	�nx��P�V'��1�oh�M�n���V�������_- �L|��y�<
\���0	i+-�y�h��X����$ۿ{�ݴ�:8��k$��2��(��ۡp�����'��7�Mc}fU�S��w�<�g�X�}�Q��9�gh<蝛�2�t���藧���{u�kRM/�̼��>�`��;���RT�����Nd����r�s$:��I��/iÈ�5n]�>�R�}�V��huM�9���7�AJdUM��P��p�o�#5�<	���l�����x����_):��o渹�ջ��a&MD�Sѻ���(@ili�d�K�#���2��b'���	�7M��]���U�)+`0&18�&��ޚ[���l��
6
tji����C���AQQk�V�F$r�u
}����97N9����������1�Њp�Ek���ύ��P���Ex2	�X!#ʞ��wN9G�W�:E�5����d_%e��}���\������.0Ĉ��m����x�ˈ�CC�_�̛x+��1���CCk�����:'�I�A_�� ��:��_��"���̾��)8]�s�(�� {�s)�͖ik�!�$�<}b��� ��Rp�Z�gG�	�G��}K�**��"�e��~U�=3t\� y��`�M�Һ�?��@�!N�Z7]W���>���5���iU��>�j[��YY~I�p�(�����RwH}}@y�$|��"!�ۻ-�J�Eکo�O��S��MM����[Z�`�l>�R,��l���8^��4�0V�����������.���
�QBup 0@��K���p���qV��cq�;����(�������-���/��=�����a)D�-�#��+���T����	z�欇�Gs�$���/<�/�������Ņ��h��}*'����v"�`
��hzYMѪ��@g,u�3d�˄^d?�7��UU���c��?����#hfd*8v�-S������?��&L����J	�u�		qE��N�O��qfF�a����N,�+�Đ��9�B�5�9���`�\�|/q׺pBl���G�@��F�)99V�?�g{xµ�>�v� �� �_ S���pWC���1P���F/�:f���J���E-.�H��!��?:R��)���g|��U5��2��~�׾�7,��5�n^=��Y�j����AI���Ώ	��#Qʠw�z��}��@(�4�S�}��퓵����P���YY��'/�̒���	����ȼ=^�+y�x �PWև�����)������c�O�ʆ����*��>~ĢD&s���/����̣o��������3�	!!CW7��F�5?��L[j\���w��zqh]����"�S������Z �; Vz�h���/K˵����Gx����Npff�:wbV��;��o(]����˫B�v|�O@�������Y�.�v(�d�+�\�}��/hs*UR�&����C�5�������q�͏�V�s���nY����C@B>z��{�j�X�� ��"jk�������a��jx�1s�}���c$߫�<�r16��OH-�/2]�����#�tY��0�̆��.i��e���	��Њl���{7�[m��%�g+;�ϛ���7v�����C�g[�K[�|��Cx:9ȯ�l���Gmk�捝���y��!/�����%Bw �q��ӝ����@�χ�b�����?~4�h����p9(
�٧�*l�+���pI�g�W\��8jC.Ѽ�i�}^������K�F|Xx��D���/_՜����$�[�'��;%���i/�濷8���d�������D�"`�^�A8�ț�I�ФK����*��#�;��C�����z�$�Rt]S05+~o�jq릁U���څ���rx[��uz�/��3?��F�o�aB���JIR�=w�����3�&8���(aeep�~���j!,�ݓP�k"�� &,s���W�׊���}E��o��y��W���S��߼<��U��ً��cf4��D�o��H*���WF���jSg���_���*��l)��]����#ʑ���_�O]�W��s���?~4�h����GÏ���M���ߎ�a�l��uX��-͎���l��̭춤�ͫi#*�5J*$׻�'���=7>}���H��]�t����r'{J��޺�YZfO�?��\ɫ�hc@�tɾ��������9�E���d����fA���߾oW�.��}Sz�_A}�?�w~���n]���z��R{ǿ��C�!?���/�Ή��:�������bZ[���a��3�v�cA�t��3y����q��?J�?�<C�r�'����E���A㖱
�D�n�/t��o~%O��=������oK�z��=���r,0ԟA�2�}�/fQ�g��x��T1�k�G�]�82</|��-����]�%0�i���}����GxS��K��R|�=@�a�uP���	1�ӵ��ߦ��
�?��n%ħ������:p�o���8zǂ���!�v���E�n����iu��(��c|�m�S-+�ݲ��	�!_����f��ㅥۺh	%�Rz�Jo�W~��WҐkX���8�c���q1�׹�����s���y��'�����M�� Ekk��`�u�}6;j�Cy�wi �*��v'�� ��P�l���{��#��<��&[�N��������P��3���ko��w������Փ\7󦾯!3��]i#ݣ���$.��mm���k�k��/�~���|K��ϯ3��v*==�5*�E�L�YX6 +G�������l.�����2g��Q8��p��V�J��ފڪC��`�������!��T�?��ҡ\�!�)Bis�N=����	VK��X���3i�l�nn�ο�ְ.@�?�-���v�=MG��@Կ��09�7  �B����d}�o6O|�VV����X�W�����9h��G��$��7���Ѷ����}8�g�0l���g��*8W�M�zQ�e
��x��ů�j����u�BHޓ?}��D���B���`���yݡ�8l���.���b�z�P�Z*�*^T@�}n�4Ag�Ƈ��q�X��3*z��ތ�Nq����&�oKуċ`����4��$,�#�V�Y��_�0����w+IF
���������Kҕj5.�c�V���"l�F����̬����L��QR�Q#e���D5
#�Ѹ�՜oU�8�l�"633����:�(1��!��fߓ���.�/��߀M�ih�W�tLɬ�ђ)sү � �P����+ ���Y��?�N���m�w��n=��9B(�Tm��Q�tt`�N+(�#���n�}�Y��!�[���������/��I�zT��q�;��9�|1o�@���ܑ�M�kdp�%����Kڋ/�#��������v6w]��0�
�z�<�)���rVwqϩG;��@M�X�5Vhh�g/��i��ykg�|� 5��p�\F*�k�"!E�
�ZsM"
�9R�W͟��oT.���"�G����1����_����j��(p}��鼶�e�l�>�g���j�| ///�r/4!G���q�s2�kB۟0����L�	x�0x���DW5g�G�MM�����誮қ��r�����c��r�a�c��'�R���6���D�z��S�������5�T��%~��}"�8�;��9��Ւ��:�Yg���#DRBiH����󳊾�8����`Q��M_��jJ0�2�Îr��_�x���a���s4�p"������W�-�5/�mu�K~�\_Jj�������P[)?]����.�uC����o3=ɕ^IB+�J��� �E|�a��TýL��hX��o�<�X�}��0o�����\�V�}o{r������?(�]�t��2í��N[c�pؕ""T�,9�kq6.p�"��3�Ш�>$��%�4�������R�<4c)zo��'��T�����x{���JJ�(5��=r�6�C�7rd����cݡ�$t��?���%�X���?h�����BG�T�g�	m����Ӱg ^M]��gGL���,�͕g@�2LM���G�y*g>���E�!�����/_�w*����=YȤȻ���N�t�WfQ:�b��R�~�$ �>�ݒ#-Wݏ�}��~Ԙ�:���959��"m&$z������J�R���W7���m!��§�.����1�h���u���qn�~���w�Έ�ώ�[�m�'?E'��o�ldK鐐�_�R4(W��{��cN���L�zJ*Ȼ�;[�UXzJ�U2�'Z%�:��?M]@�Ss �]Y�o�1Q�t�C�J�<�*זTuWo�� p�K��^��Z���XQ��(�샙�(TV�>ޝ�&d#��Ϲ�ײDt�*��3cz��?�����Vt:�$��;Q����g�ec���6������B��iR�*	mYn�Qw�8s)�[�/����%h�� 7�*�Ce��ru���M���c�.�][�qMNY�k���fh8�Hi]4�"�7#�\׬���󠬺P�u?�%����zr|̯!p�K����o�L6r���0����E����C�=��f�*Sj�o�Oy�]�B����y��;�Dғ�^��kg�B9k<n���ac	��R�05�2`I=����m=6N��8���H�]������X���n����;��L���1��`B�3W�B�x��?��H���u��`y"k3��I�����}n���s`�&K�i������A�7s�k�n
M�ȥ� 
�b�5��
<uk�R�]{�!�rH�t5��G�W�
��[�X�� ~��2Lg�y;�9�U�x��1�y���<�ј1�B����\�!j!bװ�������C[n1"��D���k�L�j��gT�c������J��A�FX_��B���JN��7�mء	�ZZ���̒㶀����7���{����r!s���h3��}��]Q���L���/D\�(涣c��:mji3Z������syM�>xN�)����N����m^o� ��E�G�<s��4�^�#M����,�W��Vv�����{n<�-�UYϴ��������Gg6ku��8�}co':lE��]c��NDo6�X6[����ԉ`�Gc3S���
y�&�Iگ!�40/���N}m���`�fc���QU�Jo}�X�n��.6�9#v�B��.�w���fN�Z����X{t������ũRݽޑ}O�gF�"��ڒ�2Q����a�訕��SkM����Ϊ�w=?�@ ��cDZzO�Q�[9�XqFޜ���6L���G2���K���C��N5?	F	3)�N|�G�C�Q��k�_6���;�`�u��_����
����5 5Pl��{�=��ru�r2����W�r�
���ɵ�1�����Rg'����5�	p��	Hd|d���1V����R�D��U��C��m��=>���t�/��W*�F&��ȩ�cK�?��1��Q��a�2�%R9�f�Qoa�P��k�tơcx�vv�y)U�p�J�)A:r��ǒ>�]��ɑ3�z�,�l�"cx X���������
� �7[�tC�n΍+kn��ￋ�pj|n��}U7q���u���p��`ܠɷ���˂Wc�@�5%�Y��H���l�����8=W %��*��g�^G�dr��g���
/]�Л�T���ɰ(b�c���4�	�߹/
#�7�	p�����ԑ��B�{��G�S�6��j�!�9P����;([�8*j�].ɔl���j������&|��P�>^WU>`B+K�R!�VW1�������-g��c}{�[1eR�z�&u��NJ��I�zh<������<�A��(kH&�OΓ���5���H�,�"�3�A�h�	%�H��1�ϊ|W
lI� �O��	��F�KB2�+��<��ɵ���Z��ե��
�\
�5����%���-N�V�����Zc����~���V��G5���v�Hb���Ȫm@v�H���L�DdI��z��cLu�$L&u�,1������܎����][�Z�
�S���E����bI�^F`� 9����!A3/��4=W�U9Z�%��OԽ6��'䈟w�;���6��L˜2�ᰈ0�zg:��q�ȝ}�lhf KD{�����^d-J�e����]Ϣ�I��A's�]A�r?!����&����t�U�P�o��CnXw9'7����r#� �� �}�g��\=(4>?um<�PU<���\���9Y�͡�l��{:��N�*E�l7 r����
0P�	ޤs�KZm�����v�Z�!A2�Z=��Ql����I!�6�fM�R�t��q�ܓ��5�EQ��2��ݜ�F���Օ\����R��b�5��}��vOS���O{���:��U!P��.�_��/�����ɝ֍��b��fT�VH�8�K�{��,��0�K>0UL�/U�
*�WQ28=�}���Imɭ1y���t���ފn72�SιL��[\��4��"��A��<��l_f�Q)�fsŝ��֩��vO]��"zg�, ��h����u^e�g�tna��ֆ+�@UQ���Q�yeР{����)����ͯJ��O���C��b�#E�M�_�O�O�E�"P��N���n!���$OO}#�*�*��(�;js����)��ݬ��uS+�|�֛?ʕx�J�<��<S���0���u���̙�!E#T������?#������Wsbk!Jd-jӔFU"7	��{�� �OPמ�p%�а<�|��<�����d-�+ܣ�;�(��.3���^�o+���]��lOj"K�`�����fN%��=�K 3��=�i�"O;D��'b҉[�_�H��DKG�o�-n�}���=koy��><<��d�^���
#��!Ϯ& %k�<`��7`�[�}��,K�����p�ii)(�1F�d~�.����������s��tu�F�öx�TB���Ok�km�´�v��p�K�u�K%���L]�^޷o_ۣGx.2��!�fF0˟���[�B�۶�I������˽R���o&*���o��vsPu�!�N�Mp��R4�i���� ih��?�8���yJ�|׷�̏{KsAV?�3��Ckv�o�V+a6I�p^��v"��u[��=�eS�Åpy�ź���,�����7�́Kp�ϳ\a�"���"#���8�b\��OY[�@�Gl2\C���>��q�w���pB�p�M��9�r]i��>3���T��=���8�Z5Y�ցWRG���a]�C�?����E���<`���͟@EԆI�ێ�}TʉH
��8x0�|]]ݛ�{�y}�F��]�����wv��p��9�)�b4����DT�9�������,�#�a~+m�H'�m��>H��Ycf�m�5�m��V1�jw���ȍ�~�:c�th>��tRi�j(ď,����)�M��E�hm���|:3N�6�Y��=\��DS)Xim}(x�Xr���!��������ǰ[QS��~��@��T�,��/��V��|1o(�)IiC�˜�}�q��%e�o
�
�ॴ?&��|,��vo�޻m�^a��� L�A:U[Y���\�z���q�3�r�н�rۯT���>W&}����!�m/W[#������_:w?� �'��?w���Dߙ=J����Sf�C���?-֪�6�3��Ƨ^B�8A*�UI��ǝ)5X3"�dY*�=�o��x���f�vG����CYW"ݞ���9���8�_~����ε1׽�5�a�7g��U�|��w�&��]v����q�Q�F|�;�_�3�ըk�UK��^��}3G.�̆�!�Ŵ30�nb�.�4S��l[U��v�cw��/��"VkWo֣�)Z/W�����
N�d6�Z2)	)�K<�3����X{ �97K;��&šKg����0^��&�
�eg ��5�=��Wx��4���h�����X�13����rL0���R�����iG�P,kH�X���l�i#,�&z�7Y�"Yn��A���T�ҝ���k˷�ƨ��#��Dn|��[��Gr~C��e�}��z��{s�R�ŔsD�蟍��vQv�HQN2g��&>�����BF1��AE�V^��Zԡ(�@��D�щJ_}N��d�J��h�{r�gl�qr��1�!�$�8��׶)�l�����gL/��S�6��I��cdR�� �<�h����'�y�=��W�BU,���B����7��k%s� �Į~���l���O���v�K@� �8��.�nZ���r�A��+I��G���>��"Z�����
R���ۃ�Cq�R曂
'�"�s����TnP�@w����8�9eiޞ�!��r���}�������T���d�Y�9^�q	0|g�p8��(�f��E�V��y��\wv��F�H����E_X�!ŋ}�3h���w�o>,|Ho����cW]��R����ցd���TT��Z�];��9��[q�0�l��ug�`ZOv^��߳�9+9����!�=�$�G�����XG���fӍu��m�����&V����7H��l�=���U.+"$_���!�d��N�:c����t�a[[�$)�1��4�%+P!M�(�Rh�����"	��ם%�А�b��ܯ�����ݰt�ﯰ��Ոz�,��7z_��DVu+����>$�iC	%�p���K~%�T�r7֛R�I�{C^l��b�����5��;j�j���e��L�����������3��н�0M����_�aIHh'�x�'�4���V�1�~��I��rx��W����rb Ѐ�!�/Μ���ǩ�|D���r1��D���yU���ג��Q���P�0�20���{'-n���Yí������2$�pC%�XQ �kɖ����ĺ9�<�4#H��}|qi'0Us��ކI:}H�md��?��{o]��$ho��PR�^\*)��3�U�	�?��S2W�8(��(NK+;w��UR�˺o�M Ū�S��=� �i��)TeR�*PY�lS��ag�Hc%�C���<�h�7x�[�7���waԣ�dy�M�b����E���E��sySu1�~�/]W��&���b��j��� L]ɂ�yO�`  ���8Y� �#cA��PD-�K�&��thUT(D�%+j흏^[���Ҥ��<w��1,�PL�]�[����5.H�XC�����7��Zs%������ �Z@WUi��^�ʺ�V�r��#�u @�'TD�� Ki�A-��+��b�v��8�K����b��{K CL�=�C�}�ۢ_�W����iNW�$
�y~� -�+myI�1��ACn�
r���k4@8�R�/lj�N�>�o|�&D�2i|�ф���	�q[�4sZ��a���_�Fs�ܢ�Eş�2˛#�d����A�H���6���-������,��{+�P*մ���o�3|ti7}�>7���*�B�C��.M��s�1 MT^��n��^LI�8(\R�,��V�EnQ�smm�t�e��ڻ��U��e�W �tu��Е<��h⎛o/X�f�"������\�4���:&ƚ���k��q���? N/�Y����-�ϖ��?Y'j�I�}���!A�Hyt�^>QI��YG�>�	G��eD2��� e���c�i;�B�T�|'�_���9e��<kȟ�\a��)�i�dT� �-�x��P���.G�2�\�l\�o����:�_֛()Ǒ
r�8z����O�c���RζE=�#�hB�����a�r9e�r�M�Ų�I=�d~H\�z��,7q��p������o��VQ���+.
�<�q!�'�`Ώ?4o#�HYov�װ�~{�}�!�?	<�e���Z�
��bZ��Vɨ�b��,$s1���G�5=��G	�K���� g(~+��*���HX�����������o��
^碋2��~�Z�K�*��Z�geĜ��ȷ�^��2�����x�y��	���M�^�����w\0{&�dGQ;;�'i�Qr�2�j#CnR�F�E�ސ��_n���s��a7��d���w㘄��g�S�\O��H}ڸf��>�~6�,���-{����D#6*�T�:r�[Q`��'B��$�f�����}�u�G3��=�n�mJ~�f	�C0�}t�%m�,ގ�y
��C���Vgn�1�Q ��bh�>���d�nv"_Ty���j�4��N�y�g�k�?�?�Z����sPz����E��,����N�kݲЏ���r
�ė��Y�^��-B�>��0�{s�ya��#-�z|�:�I;Q?�v�'x�ި�B��c�	������ͱ�Q��k�4����/�c -�~f*��7/'�;MbtR`Zv���xs� ��z��r���1ݢ[b��+5�ۂ�Wŭ=;3�'g����H��!���>�#�� ix�����-'�P`25�K�%�q��K�`�C^.rR֡q~����}o>���ܵ�1^kw/NA_ 7�~k�X`Pe����x�ߗ+��3TB\��l��7V�1���l��e����9�n�n��TXܵ1�I�4p�!�-��b�"M.и�H<sK_"g���b�!��d�T	E9�������N���g�eO~��SU��o$�L�\h����yM��A����!p���X��������g- �*�h�$�@	@�Bi���ғ�'
�
^V�3P�Q5���0+Uh���j��߼�_��+�T|#��琾�9�w�Nă]��3��i��e�g`�3NL\�;�԰���X)�c�����m}u����I����U��&��9?����[׺s�`�xw�C�,mk���A4	�y����F�g1�D.=휵�0��.�l�'G��[G���C�I$�[�,*��K�W1@��'��J�0z8샭rB$�Prh}"T!@T�Ȧ�����v4��C9k3-u1@L��п�rQ���M���BT�A�����V?����Z�@@���_��O19]'w\�]s�����
��`�e��Hv���"�ՐOTy]��s*�26D���9��2����*�/�Ӽ�n�N����k�k��H��]��L�?���!s"8T���b.c�N� ���G��-���h����U��R(4�p����6�&���Z�7��Ȼ�.K��� ?��\�]�Y��8hY����`ň���Z\����)��o��-�9���: �0V􁄮��B@[f�U��`�|�����e�5��������\?�bt��q
�D��29��s�ff���&�͕��a+��Ha�k�?���/t����j[Pl��D/z-´p�u$��D����F��a�<᝶u1н� �����t�iL�8��o�Få�6����@VJ�����@�h�6������F�bG!G�K�{�<A��tvY^J���\_���Ѥ)�.�gk\/.�=�}����$|P�y�o\�Z��bX�P�p S`iz����c��$�שּ;�_���uĪ�x�2\[Hn�/zuH����dt6��ױ����l9(��K����^�X]��z�*A������T�K���Br��3`,�q �U�!I���٭�ut��C��ZYjy"*[
}C�A�9S���P���5��k�����؃��M�x��G�aS֋/L)�����Wcd��;A�=B��-�����/�u��T��ľ�	�K� z�T(�CB^�Pvj��D�]�|P����-e���+Y�WԴ�0�r�^�W~��IBw�|I ���{��!0vߖ3L�����Ҷ1KB0�]�4�N�ݴ5I~�:�-��X&���@�w��v�O���D+4�<`9��՝���h{�Z�'�!#�~��W#�W�`0��|�6��^�x2�2�j(7Y1
�S�9�dMv�6��Z��3�w�6�q��7�ʠ��U~�F�(`��(wWN��6#:���<A��B��
�K�Ǐ��h}�27�m��(���A!t�����שA
��^������򓗁1b���q�]���o~�x��z��p���#�g���/饣"s��W�vˈ���76�9L$`cB#}%~G���O�]��ut�P�-�L��0tl6��ռP�>!CGbC߱��Gs�E�Vr!2W�!: E�M��nq:���/�6͘����лhR��i��7��t�U���Ъ�����Y������%�[B�u�����»BP �:crR;VIn��p�q�����:?��/�'Tr�������ρ��+�*�/O�j�^�
���38>H�)�t=�D�'Ǭs}h����ڎ��U�/yy.KD�c��zy�F@P|nX����Y��[�qc�0 ,�%�&�� �c�q��5���%tJ�� ��l`��~O�2	�F�T��.�D��l1BƵ��r��Z��{������v��/�t�?ՔMN�Vn3X��Է��)��J��N�bRn��T���4�%�2E3�r�%�#�-�p�ܐ$c9������g�߼��k�^����1Z,���#
���֒� �`@��Br,�?	�C���P'��;'���`0ԸWz��x0 P���zj�H���H�)��Bq�?�;<��]"�N�U��0�[ׄ���
'~�o00���.�P��@&ȔH���]��2�ob�?Moӳyi
��?�k�V,����f������vaZS�Jч�C�� ���v�����헾z\�R��uC&�����ј2\쳣��� �~�n�S���?b��OY�|�}�攳�3���T�+=ZY��ꪂf��6;���{^,ڼ���Q��:�R#�h�$X�.�yM_��5�}��*MH�
�E��T�+��� `�tx�f�;>>44��S7�*3x���w�	\mj��\��gձ�iZ�o.�6D�����q�O��Uؠ �rB���
�ڊŨ�%� ��?�W	x ��K�\G�4���J#L��A*�{��߬8��O�mV'��O��"A}5�a�������Ձ���i)��zr+�$�!�M��t�{G�pP��yН,���a˲ngK��8ie�%�Ե9�/��(Ywar�DR5g��iM��= ;hki��;�4g���i.(�9$m�i�n�'Za*V���~Ϭ��E��<9Gx�SzČ#T��?���f:�X�;��@���+V�i�$�i7
���{�I'^J-{=�U(�[��ΐM��Q#���ۤe�Zęt�7 Ά$�&%�>��~����w��mb�P�e�d0bc���R)��&��3q�%
q�w��0�\���	~��w@��#��A]p�:�����ȏ��ҹ�e���kZ�i�<�v?�0����"���tck @v�w�M�5�Zi;C���L�����ע �^v쉖�5�B0�-�� ��r�z��nԡ��P���H<��8�8SP���Wf}m���5��r-���e�&@���Z�%F%�QQ��E�1��H�
H���~��-���#9]��tp��x�"]WU�Ye8_��{�]J.��%]Z�7L�
�I�xQ�82}": H�*_vq�3�V����;���N�N��5�X)3-�l���b!S���cAM,�?R�����^���Ǉ����*�����/��efɿ�7�p�
��J/&�H#+>^�׊~�|�j|��oo��?���=�����]6��x'���Z�Q'h�}��$Tj}?�� [���K��.�f��]bO3�K��������)�NOΣsL-���a��>?�XFp����K�����n�ׁ�_	 �7#��Rg�l�=��ѡXj#>�M��T�Kz��FIp�K�C5���F��~�B�ĳ���9��d�`�ӻE|�o�[�.�>���Lw@y�< ��	�r#%��nR�@61��m߃�S��0��X�fs+����W�F�n�sW�U����CD�%TB�
�M�
�M2��V�ع�����_dYN ��GԵF�s��z:cի�}T4��#x=9�@�Q<T�����T���67G��RGҏ�$	v��'��(��r��Ei���;Z#�ZG�.��`����I��L���]9"`މv,$�5v*p&�>�E�p @ܻG�P:v��5zPy�6|9�}P6����l��������yDb�C������ӫw焢�!{��r˾wwʄ�bL�g�d��SLAhw��j���N^��b�L�J�(~)�%���G�F��
o�3 � �$�]<LH,7m����\n�='�S�&�A��Gn[32sN�$�����(C�2���o��᱂|Ik���ݽ�������5aՇ+U�QF�n度���b2*Ʃ4f�n��i#dJ�|U
�
�#O�ͧ�k�1Y��U�"�u/�O-M�c�p�j�f��W��/�̭�.����C�fF�d�ڙ:"��SŲaK8�JDL��� @�#3e�&��J��P�-�CwnoC�HX,ۛ���{+��_%TɵѰ���x�,�	dKj��S�묃�sj�w<3�)J�=����� �	�B��ڤF�ķ��T}��������pb	���C�K�����I���{����F	�0�+���S��L��_a������B��ZU93���t�׈�x����!�Y���n��z��	�P�$m����.i�Z�#H�7́Z����z��4�h����Uְ��>�ܛ��G9O��f�[	���|f�?�oi��8x�Ax��'�ܵ;o��xUr {pA0���^��\zA�9?�P�EWI������3���V�rṳi����{.U�T���(n�7���AiǇI����p�d;z���ƒ�Ę��^M1�ׂk5����G�q����3�vd�[���|�U�1ydߗ�{�ۓ���Q���>�.�8��;���!j��?��ͩg�����l��Y7o�.�O�-�-,�vT�^t=���ʆ�'L�k.��bߖ��vR;$�m�Q�)��:s�<�F��D$�um���e���ah�~�����I���s�K����F��>�9��f�t�i�w�"u~a�5�Dby>6�]�N��?�n#�o)t?�޺҉ko�(���C������ ��xG�����Uks2+�@)u 4+ɘ#hb�۹3P?Å��י��V��	Q�~B ��S�_�)�%A��nS}�4�&��ҟ��W_��O�rpY�uvG���i�c����spt#��?�F�tg͈٘[{��7X�������g+#�J��r�� ���7�a���܄�=��ʬ-��W&�I��'�OԺN[��t��f�|�#�C��V�a��D���y�����q��/� ��<�2N�� Y*9��ħR���k�w�����/&,�	e�.��b��$������4I�M~_���߆˴9��(Ō�|!lHͲ�%����ߍ\<����� ��3Z5=
25-���OX䞤H-a��FF��	s/�0��feAK��䘼�ND����k��7ķ�7]2����'�� ���ƥ؅�Cʵ8�[Md��&Y�j�09�+ȝ����>G��
�Z��#5�������%��u�!��z3�U�-c��a����q�l��<���P�G�f��pr������4T]�����uP#M�)�6���y߱����Wiݷu��S�ع�����Z���Pt��:���i�(�x�4-C�s':��&��^���� �狣���CU{)>�Ñ�G麃���#���Ҟn��Uq`�g���Z>�#� v�kF)S;N�@��t��ĶN,���i���8�w����(�a
fz�����{�6���MQRZ�I�����{N�b�ZNH����gL��b2FW�+�=�P�ll�SV�m�$7F'�HwJFghK�_K�Q�a�&\��q�T��9Ze<���cz]Le۸�3���8\�"C�P0(��+��8:}L�]�<�|����' �C���VJf]�dV;oi�,}K˶Mf�D�����Ǵ���C ���1+�����C�ᓒJ��[1���6kKڝ,y[)r�z�.j6gL#�H��wU�ş�Y�ub @x�, �Lېd��X��rn��%���R@*͐A	�����4,�\F56[�S ~�͋� ���qj��K̘;y�|6P0@�.e�����vʊm�-�*X�I%�w���|ko�:c�u�S��#V��6���`�a��7��}@�7rX�Tq��{p$�>9ib"u4T��F{)V������W6�6�1�g��~s��Fz�C�*>�X2eg�B�Dm�(�Ȭ6c;��J���:\%�0� ��;�Ky�����ɦq�2젮a�@����6_�(��s<ξ�/��(��t�G�4���/�%����_���P�����'���$�A��t��]\��Q���u
_v��]��Lų���D��&�K	�#m Յbc}ij�QL�-<{`��g�!�ߟ!�=��_�APIZ���L4�|� ��A���dAA
{� �ߚ��x��p��H�W�����)<a^je�l�2z���>4��~a���?#�j�/�C�1y?����C#�KWZ5��h�v�9<���H�q�]��ڛ�]��R��#7*��5XI��㒁�?��RA9��y�L��l�i2s�e�3�P�5HoX㻆�VcT�hN��_����Gwb�i:�o�ji�����o��/�K�<v��D��Fp���+��I����X��	�K�w9�A�)��C�x{��(�o��yfĴ�eD0r�ߠ+���q<��}���e�����t��%!�fs>	�s�6��B�Z�E<�d�0�(\�C:�V����f�f��B��sM1auֈ�YU�J--�5M�n�Fs�j�$R����p|������?�CP�[j��L������Z���?k���']������d���<+�!gO�<˜��p?)�ۍ���g(C������}+�H'�U�K��8I�+������r���k{�R���%M�� Z�3����T�(��iH���30����q�x]�ج%�������^
�$��`����K�,��<��zE���B��,��Ԕ$�;fiM,3�U�4�߇��d1����I����"�v�J�>��^���
�Y$^�4�W��?�<��0l��~ۇ������.�����W�4�,x��r@��8��[�8 ֐�0�h���m�q�h�K�zp��mw�󣭌	�)�ڝt�w�k�"�*�*� M�5���-ՏR{�FC�ɝ�h��ڏK���HsN����2��p�T<�<����iz��߳0��6��9�����+�yӥ��RU�<����~DU�'�3Vz\le��ӈ��9�����[v:��h��z�=#ڨ��U ���m^�!�)z�	]؄Ƙ?���H�Tܞ���V�k�6	�q܂
״�T"�<�����e4߂Koȹ(�4h�5��_x�8��L{T�j��l��L�����`�47G�M�$K��f�b#�t�H�c|�LC�����o�S��)�5�75ei+�&��\9a��H��։�/5&')]�4��I��4�/G??^x����FNz��O#y)nV�<V�r���m߬!��D]xiR�3]��{7�3{�����A8ho��=?�`1�G�=@[.�ʜ��}�����#$*��	�&��{A�f<���PK   *��X�����   �!  /   images/4b131f3d-bb43-41b7-a007-3fb3641e8d39.pngmyg@SM�v�&(��EE@B�*�(��ޫ�ޤ�h#M:�""��  ���^����N�?�������svgg�yfvgO4L[����USU��.��GW(�����#w�jAA�
��S[
�M�j���I�KӎlA �5E�AP��T�;����ʆ�#8�x%�A�w�Q���6�r�+/��K�^)�C#����¸T͠ד���|�3�<,��,N!K�CW�'����ǣ#��v���-�嬆J�X攬����6ϭ�n�~N�-'�"N�T���c_0��	����|�����E���}�{lW�P�e���Ѥj��K�x�mĭ۷���t��7�}��(�#����� �!\58�8u�/��'.�L8�X�O��
r�g���,�C�!?���t�(���͉@^�7v���xA�(]��l,0ɰ�d�ge�b<\�$V'p\�������Ok(������[��4^I��G��|p�n����g��UV2�3a�8��DD
�J�M�?dt����N�%�L����j�(5�QM�>^��\T'�����&-�b!�MR�j}��^��Sc#��t	?�	�d����t8Y�^Ⓦw�B�ݭ<lְ�30}@��\���>~ʘ��Ӊs�CNT�K���>�y�^v�����Mb�0K�
�&���|�j��s��9<h��"/Z\�dOs���Z=�FҴ>���iV��
k̍�˝�b���Ff�䜅�TX����P��:ϫ}p7�����Ժ�<A^�i�@�/A��HՓ�"�������� ����q���]�QS�w����Ȍ�	�/�[�3�״�����a͹`3�$W�ayP��i�vwL?�d�����R�e]�Zʻ�v�⩍�7�_�G�G-N�c~9�6KYpD��U�4�_�]��g�+��.�D�,6��Ȩ���'yE�<%�"4���_��/h�-;��:v��ctR^��cUJ8��tBc)�� �Y�h�dǙ8���`{�Q/���se�c��~�a���B#��=����x-����$��Evz���j���S��@Ye?'T0��>cd}�s�dl�c� �e3MC�h�v?'�\��)&-m~�\�&�eģA&�i(��RG-a���_քck�(I�^
���4,��@�XǾ��O�oia�-	�zy�����*%S"�mn�&Z^��+���H�v���`'W��|��0AG�܇����#�2|r��K�.9�����Xp����'��դ��ז��>WL��B��Z����z�w�>�����-�u.�6�`KT��\�-(<*2��r�����5q�vR����pxd8�#=?T�`�c��'R�K��՚#�(�=z�%HjĚQ�J�cV��ޅ1{z�GIԓ-�*��zx;\K9S�ZE&4ť	�m���#R��o����^߈㓧�W'����uА��+R��v]D�w��[�@���^��[�%!��W���DKK{?E���V
J�eq �ah"6 D���)�j�ܖyK��Oܺ��Z�`F���&O$�W���a7]i��o��VVF'aV? �1H�N���8<�GoD�S����T�ƙ���]���k�|Nzf�}��|��1?j$�C>�æ�����mwt`�2y���3���۳�����m'l�����?M��v�Za][A�s�N����d<��<?/��C�{�&fdm�����	������5��>�L6�l��=���rR�'�9��sS��'���h(&8�8�r�V���1Ԝ��&���:��Ǔk��IGc���0+B���z_2����MR�	n�AZ|h����e+Q��V��P@@ �� N������F�4�����:G��<�?;;�ܺu��+**jdyc��tg�b�s�t��b)y�r�/ԛ)]l� `�-��p�~��4���W(�P=��B&���W��>q�9({
���joy���,%�3_>^�dV��;��8�'�K���gQA����єo�r��T��jU���k{G#�Z��C#5����͇u�eؖ�+��o�T��v)�_l@:�}ɣ���v�_xBe~��(-%����4�&&'W`���с}M�v�BGQ��UD���i�S�sLIjj��U����k�Z뿠W嫟䠁�k��OKO�Q����l�,�]e<F�n[{��0�}u7���W�#1}���yx=DBJ����<�d�&V�,������-p�g+�xvk�k�'��ƫ�:!�{� �+��;EОԄ�P�����^����~hqS�� � ���'�C�S�'�4�~hWsQ���j��#���#�����˾)F<���j:�u�*>r�8����7T���/36�T]kC�SW��{���AS^*��ή��Lp�� c�2��zJq�-mC�צý���s�jw~�������R�u��W2�(�%�l��--�qE[M��q	;c}�Q<��T����{À���v,Ș�ۖ�0mE65�h�"c.�n����%�|�v~8Y�w�^Iׄ��F?3bv��j��OPv��݋�͒�����P^۳gLw���4��qק�YY����[#T��������=���;:��JT�ɥ@��Iu-��D�]��7$mے[�t޲'Ӳ��oa�P���,��|��>�F|�� ��;{���<Ԫ��L��̂�4T�@�/0��ZJ�T�j��˚��Uq��f��2�=�D8d6�yx7��{ݨ-���W�:"��N�r1��INVH��*���%s���en^{U9�����u�����
�G��<ߚ,�M�R��S(�!�3�6��u�7�ߑ�Ui�='6J3K��Gko�?kXI�m1��	3����m�{%%i��nw��Q�Bx�QKj[+��4O1��N7��-��b���	)#/�^��#�%�r6�:64�rs���}�95k��/�Z�Ԥ��wf�dJ�\\�ƚ5��5T!1_95�=Bוeu( C�[a,��&�F���ɽX/g�Ҹ���*$��
e��rCbg K��+E���uڦ�����4`�]������jz�zU�vZ�YKY�c���U��o�z6�Z>� �v��+++L
�g����ɕ5�<^�
}$W48"�Jt�V�P�4�L��0��~�~�}�̪��Z�c6݊� �� ���͡��|ھ���Px��X�b��V�H�F!L����b��G����ngy��M�{{��O䀝�_jZ�^Y��6-=J�<�xfMXf��`��5�-苼�i�߿��H�/!+��H��V�6g�q����?���6�z��5w��WG�[Ͱƣ�M)�^�%�s�#1�	�ݦ�E��=h��U�m.( 箋)58ѕ�]ӽ�H���sd��=ճ�6s��Sd��{j�7��Oi�k�i��?����yR���qL	F�<
*2�	��0ٲ�'ڂ&{J�<�@ �X. I��@
��%|��^�v�RsOG=��s�@RTG.�����۳l_��nt_@D׷��a��=)%,d$�E,�SS����V;iƺ�M�|	K����e�����=n����j��!&�ݮ���A���ͷ�-u|_�I������R���Nj�C�ޥW�e��`8��8�HF[9z����i���[���@�<7��lj�f2�r��#�����`�+B梯��������:�ϊ�y���OB����:� �B�g�_��^�f�z�̓Lʦ�o1��ucc� �VC��.�*��r����𘏑�SR�t[m0��J���S��m����|:u�2��E���	�o�8oM:����t-T5�Xe�b��Q���Qt����~:��=}pS$�?�ꑾ�he�T~�&h�w����������?M��]7���֑'�si��Gp`K{��x�I�����BTW�Sp}�Ø讕��eJ`��zժE�L��GG��D�v��l�[�LY���8�V�����K.�[D)�l=�5�.�c���^�Α�s�����~��lj�z�`��E@L����g��oN˖�`�m�����[0����r��d�� ��D�f�Xe�
z�۵gU��G�!d��w=�����2\2��y�f0�&�/�̥�\�W���E��W�[h�1|@Ǵ��D��G��<�OH3S��?��̖4�VL��9T�@�ͮ|�E�}����}<����`�'�2�͒d�.e�=�m��"W��2
,f_cb�}�h�ε��G���n �	����q�I'��-������‭F�wL%��f�=�	`bC���^F�Tf��!�LO�,�j��puqQ���+���@����>�n1��'�O�\Q� �;��c�L����I�Q2�߸��6z�c�Ziǂ�
��|�kM���zkZ<Zt�od!�N��T�LKQY�Aw1����ӽ��	�
W���g�ڽ���V����h:�CtH�����P���W;�AS�ΐ�Ō7�]�pI���5$��YyLT[��rrR7D6�f��A�~>�do�i<��`C��5u���>�kA'��>:�4��*����m {���τ�N�X�<��a��9�S���S���[@�p��HyR�?�3�AO�U���}��k����2a��g�R�g�q>�z+�{I	�S��F���e��a;�ء!e�r����ꃒ3	-�ځ�gV��gc�2�Y!�j�[;��R�d�� �J�:�cT�S�Uz���G�����-�u!��	̋0'�Ѕ8�Ȟ���g���7��2A<�_�K�F�^������ކA�#<?+h�E�6�ج��ĸ��Q߬����l;H�f�t�T6"c%�ܰ�>�f��N�s�.5B.�m� Mi+4�u��@��`,�;����Ճ�e�g�G�o�'*J�ݑ�U�=�<��?��Z�	j�$��os����F-.A���J���/�;ܺ}$���t���A��6uL��pn�����i�b�w�C�]�o�E���: ��!Ic(K"��~Z^g�'J}��#o����""!Q���;]�ٳ~�֥���w�hٔ׭i��3|�0�[
���g��Myi��Bx����/M}�-����&%�s�F`Dm���M�l�k�٫�g���$w���犂�dl�Zū|���c����J�z�����W�I0ԗ�lW�̡¾sHRˡ�gD%{���ყ��KjZ��A}Mh�y�6�m�*��G݊��>�&[�x�.���V5ǆ���ӞgYƬ~n��þ����@��ЀQ#?)Q���W������?�C�*w��+>"��iT[��&r�$��q�k쵷���>XmR���-&s�����H��j���GBg!�S	+G*.ldK�P刏1��N���\k�Ā���<�AhI�|����QGW���gr�Jv�@a{��Mv���I!NLӫ �|�
q��W��^�ݭ�b����Fݥ5-h��_E݆AO�E)�S�q.OR��a�wC.H��L�0@�LF�h	����#ԹX���ܩ�7�7�+�kשZ�[��z����)���U��߯�@�euypnU�4F@r�c�:�q
	b���&V�$��_�j�-^�Z�P�k��}�ǆ�JU҂��y|��1�t̪Kau��dJLLT�v���Xh����s06t��z�u�|i�ALȾ������YC�u��?1���m�2y��*�<Wf��1![���>f��I)���Wnh�o���s����s��(3�'�0ClD{���0�Aj_�z1#�S�5��9��b�>=��{��v�-淉�}�ݻ�z�/�Y-����ӟ.�Rm���ә:'���;����'�5����>������m&�ʼ���0�̐����l�|
 ��Kr.�f��ؘ���﷧�,�!{��f�*,����k#�wA>d�;i?�S�o�������j�+�|�h.�S\1#\�Z�>:���[�}^�p�P�^�B�w96t\aqX���8��iKLC����΅�?紣�����{y(�seű�����󛣂�G1UmB��G�?���̚���=�')�EfW'Vm-�5�T`��
Y="�nii��k����b��\��5݉�*l{Qӄ����41���q��Ϡ6���[ob[�b[o��ZUz<s��_��樏a�,t�y{t��q��5��Qii�?�V��y�Fk��l�N����ni���f	C���1TA-}UK��7�h��8q��9����i���'xLD"�GަO�
�6oJ�k�L� Jz3$K>�]��%�E�V�l��8D[�9W�5y����-�u�u��+����p�����b�}����͝�R顂�ۦg�����K��K�T�\���7� ��g�p��1�#*����4�3�.��x�3�_�DD��򓭦��W��*n����#��M;_ƿ��U9t�f����9T-���>Xt�����E�sq�ݭڄ��7!&f8���bn(}�#���M1�g���L��O�t�ſ�]6�r�X������(��o��?v�X�n���/c?��.d�<E���Ƨw~�g:B}�������ܖ!kn�0d��,���0�.��@��esN��uF�����PͿ[���;W��%�/R-v��˽_�?<~����{$^��-����������6i��D�W����a�T�~�C��c��1���m���~5�6�_�o�͚� t�F��1bQi���y���>�N<:U��hxOǛΈ쵑H3�f�ٓ��gXGUa+o���)+�e�=D�_�ws~�(���ȇͭ^���!����M��>����Q!N������ �"�*����F�sl���y�Zvԯ��W1�nR�d�_)��6� �Mu��WyJ�Փ[]\K��I�Ei��f	Oa�L^}�3�y�l�Ĕ}I��Ѽ�E�ʬtx����?��;H����^~i��Z]���=�H5ʏZ�E|��(����T{�֑�[��!��
���VH�1�
7���� ڤ́��;^%��6�/f����|<�iuZ=^[XE��>V�ɍ�"݀��7��EwIb�1mO�����K h����:�5i��9^�E�:���߀�x4�m@�9����tL#H��f����~#�$�w��t�suph_�2گ1�I�c]��\L$ �5k�N�A�f 3"��sH�dpR�W�^h5�H�$�����������*�v;kv'`r:�����c��$abH�2-�x��x�"M�|>I�h_wÀ�G�q���E6��h5���v�����w/�������xRhp�$�����I���WVV���fw S;:;˥�����EZ2݂�"���RgL[忟.�Iz+�9�aL3��H�Њp�,�;��ɯw���O@��߆��9��NX��r��7zE>a�'K��b����:8+.abL*"$��k�^�E�W�/�<�&�zʀ��=֒!X/��c�'��rIgU�u��\���������$���Թ�Hl�Cs.:��D1h� `���x�PN���׆�����SQ��
�%��t��t1����7�z��v;廁��bL��R)�P�Mzdp؟�oS��EwG^�]��}���D.�C��R��G�=R�z�T#�)���iy{�L���1���Ec ���L���$�M�F�*XQ�%�Q���@W�Тq�jCx�t�I�"�P��\�$�?*���z2�#I��B]��E��t�%�t
����D~��h�8�Ӏ�E(��)�d�2�0UA��ܙR%W@/��хCC���0�C��dL�]��'Z��DF�R�(��-
���"�1�> е[@9���	�%E��N*�:�T��O���o�*����Ƀ��J�i��Ѫ?
Hv1�#<�C~Z�q��
�_��@
���r�G��NH��
��$�H&QXI'�|��l���M�!J��������@�j������V���_~��&7�\h��FO�#��Ph~+{�<FT(X���`�6��y�p K�s.�l��u�>��W}�\0����g�	�!y#�֍����z�u���@q�1r.�'G����K ><��T�U���#�!�-PT���n7g?!-�G�+z<�����m��[�L��G;�qsuN�8:��TW��\�,r�2c�"�F���5��˖�Ӑ��O�>n�r��%��t�K;�כ�:/��eh�<6/�^yIz���	��+�HY��¤@���΍K �.����R�A+C��4�+E^d\ɋ@�+��u����,Ћ|T�$e��;$6��S����j)#^u=�"���NE��O�`���+�nM�zT�I]<�)i+~}b��PK   ۍ�XS�ѝ�  ��  /   images/642b7e82-22f3-4f40-989c-bd067878f1b6.png�|�?����:*��]t���TӉF�۱[D�-���d�4��w��!Cw5r�Rc�RVSİ�H,Ɔ�f�m����~~�����^���m��z�_����z>�]�?�{8���U��������ƮY�];���y�w�5����Z�|mԹKH����ϲ�P���[c���\@���F�����F�!���"������~w:�����W^c�J�P~��.�ݪ॓�Nt���OMǱ[���{t������NvF�ܶ�|��r�O���\Y=�n�y��'ZN�5��r{����b[������4^E��˩s_j�}�Q��O=�lů>���0�=�X�b�2@������w��w�V�
j�N����L���##�PB4�i�G��5�nw��j�U�;�h�9��_�UwJ����X(nU5�%���+� y�����U�O�#9�ff����ϕQbA�x��2P}E����F����8���r���曙I�R��kѶff���^�i�)�v��Cœ�:Yr1R_�B�X���uZ�n��,�\f�k��L~���߆O��7��o�m`N���,�I�rA��=xq�d}E�!k$�G.���UiiDA�Vk��H�̮�2��ĜP���� ��I�vvv,r]]Jaa��i����	�ǁ@RI�+��� o�����#��l���cp7�p~��D`l{17S҉��-�!0�˄ؿ0�iC�f��ӎo"��0��f������Y^��iܴ~s���)xd����-�ûxdF���d�̮�����֤"#�W_���q��Ĉ��)�8B=μ�"�*���YD(����������։��B���xL�%?�[j�Æ�
�S-"����>C������L�P*��Ԇ���RY�]�3L12' ����?���@��do�BX(����p"��_��!��[������~h[E.+��5!KD�#��;�F2["�����(U'23:qi�=��]�b�Ǧ`�f��M��,���������� Tӳ��������i�����0z]\�/4�8n�V�A�=F1�,葬�?�x�멁���*�Oy�D��'��~�C��ѿ<�M8�~{b�_s�)���s�Ć/�S%(h�(p��[�3�KQ�8�B"`-�?LY�4|��me�5�)��b"�H1'�
�=�|� �
���9���g�1̄ ��e��N4^�*�M�Dq{��mE	8�aJ��-TP��d�U�/J�x�3A����q���e�w��	C���9i���P`�pؠ�/�X0\�e6S�e�y����&}{'o���k����@�����	��J����o��e
�I���C��L;jĎ8�\�� G� �0L��B`#�`ǹO;3�;�M�Ỵ�zE88�̇愷 <�Y(��E���c�6}}�\}�}33B����^�p�j��f��z0��x��9��^h8��m7bZ(���T삂""�*���&r�AC8��� �C`��)��?k���wgi�}�%
L�RF8�̮���B`���|hOc�v!��,z������8��ل�ؠ!��H��M��!�J ܪ�@]i6��.NXۅ��U|[�i-u� @5�()�Ď��0��P��\2�>ܵ�k��[�1	�&6����W�qJ��	���Ԥ��>j��U�)��(�t
1��3�l�7'X@Y�|$֎sՅR���#�����5(�#ip�me?���v\S�P���&;}��� 
��Be��w�BeÖ:z�N�z_|��%��̞{��Ѩ��_��hMz���X|����A |��e���$�Q#ge��AQ��5kA{�14�BY�[���R@7��c����J�f�.��d�?�b?>ot�5:~�8����݃x�,l�d�����{Uv�?0���F�8@#�ğ.�E2 	7��/>���G������|�>W���\����^�K�ړ�y�:�6�x$P±��_�t[Du�P׭�z��l���N�@�5�,T�:�IBAeg]&$�XtAd���AP]�	��u��=,��*�	�y�a�:@)����4��R�8����eN�e�.-���W	�_7�<j*�.r���.��0� �F}]1YA����Cv}>˛� �ě.f��<�M񳟳��K�M��H
`'Ȝ�J!��j.ݙ���Q��4����r�c�Z��2���^Hd�|�� sb��z�(l/��h���Q݄N-���ǝ�������L��S����p� �S��Z�N�[���E��:GtAM�6�I�7���}�U4F���z������k�C 10l@>g�����E��}7����w$�i��ٍ�r#��m����#} �6gO��LR��q�xߵͪ�ќu�?i���;�bPOR�I<Y��l��[��UW��id2K�1����Eq�~g*�����L ��"3��A&��a����`\�|��lp�\n��\n#�q���o9X�l��Ъ�?�ʔ
�z&o
H�lZ�=/R<�21�ǆ���� �p= o���+��b�.�;;�K��x���>����8퇖��qma^@φ�2�ޛ�p��"	�Bu�U���3�������!�'X)i��h�򽥎��y���v#����D��;��NQ���w3��@3��s�X[�""Ϊ݆��z6<<��+�:֩�V���I+�
=��龞���������J!h[#�d���� "E�'23)�����Y@7��dC��#��M� ���-��Q.�Ĭ�^&b~�%���Yi� u�� |T��RI	+��)T,kV��Iť����h��uo����Y��˪�.�"t@Q	K�-�]�0'�>`��dv0[e�fY}* 9��)S�\�
�)��tZ6ax�EH�``&_��������G&7�A��h�i���L:������@��G0v��I��*�|Es2+�\�2�L�s��@`!�����?���R?��zs��m���BlW,	����kn>M�>��^����1;���޼4z@4�]&�r,|�
4]�&gܒ��iǁ����?���w�de���r�eQ�#��Ơ�� ws�A�A�1��{�����ތ�H�s鈤� ��)��*S�@HkSf"��sRQ���I�&B�a���zCpz�[����=M��ׯ�s�z������1^��Z	�l@u��g�1�W%��N�31��Of�~��)Q�=�a^�Uis4�0�{�Q�\����̄�f�Pd��X]��PF.,q�jc����Q����(o!��<�ҍ�ׯ��Rj��g����ج�[��x�=9���
�*����ig6+U(=�ad�/�kN���}S0�R�`wFգ�b��^.�L�5�U��Gy�i-1�bu��\�S/�D��]@V�A���7਍=�B���?�����A\���|�ȱ����[1$��m��f�aÜ�I�٩E_`?nN�9�Ց�h���b'�R�k j��0��lu�B\o=�J]*�l�w%��v�s�q*?��3@)��h�N��e�G1�����'����S8y��,O9ᚯ���0@�B�%HI.ո�R�0T{�*��DJS��X�5����.j%@o��pN}��{y}�t�s�o�gi�C��GO�Q��d9�<����!#�F����������؇OE��4�B0nd|����3�.E��9��A�@9�3�:���NK�9�����t��:����_:�W��~Lb�f[2Eb��e���X����m�>vG�:�Γ�2~�w��Ͷ|�ko�A%?ӂmf����U_���2I���-����}�7~yfUf(���q4�@]���=�V0m:������x��|7lЏLgZHIҷŅ&2����S�'v�E�i�/�����0����岴s6דћ O]�QҺ����9����Y(��9Ƒ#�==r�`���2���`��?��g?l��Eq����X&]S/�6�o������z@^��T����?�Ť�bF�Y�L@���5�|\�W����O�o���T�����?��07S�7���S�';�����h	��X`���/���B�Q��L������E��Ft񆼅Vk�o��BbcM*�6��A����׆|j#��8V��hI��3uf�gPh�\@�I9D��%UH'�%�!�fEX�+���^Y��)k�S,!�T�D��J�@����^�(��������oD��i?!Ɔ�(B2�(B4 �Z����͏�q	�z-Ļ~E\U�Iv7��{�����
�$��߆w��A�T�z�����i�3��c-CV[���z�}<(�m# @ל����l�.3���[������іyU]�g�\���&UD�:-0<�@x	�Ƿѽ�	���*�Ҏ^!�k#�t�jiZ���J2_f����@�Y�K�R�_L��fRM�Â;�hާF�	 jt���v���F�3��hf�6�u�����T�h�~E���0�,�>�ʕ�Z�� 0�/�W�"S�l�q�Q~��vO����tΜ�f#�˸����������� ��v���a��m��6���) �GF!�[c�)~��ॖN�h�'a@C�,B�NˌS�k���S�N��m������o<!v����w��\'��j's	�a���͚R�>I�X3U���>�l����1�$��}h�Ǖ]��뤿�A��a���ܻ@��.WD{B������2�2�CUlJC�����ľ�^�
[UB��!���I��y�����DA�n�%��䪔)$~��� �mw�D�-W�͜����⦧��3�\�T*����<JY��M�%
If�OF�mQ�@��Gg�?Q�����B	���"��A�=`j�@��"��w���!���S���Z��(���q�w/�&
����h"-/�Vy�Hi[X4@�X�������N�`�@� p��(8��f��#�m�������3NN.�;	5P�����Ӫү�^�I��������@C�P�?Ӽ�לܬ���C���;.������O�]	�~��C���]!�?�l�WT�.�@_���ؙ��u+ϧ�k7��݁�q&��vAm�'��������ێ�v�k�ţsII�vN�_�q8��b�rY�����R7+�=1'Pc���f�b�ϐ�<���6�D�Q���݆K%��v4��t�W���=}˜pH�Yii�H�B�7K���/<��E?��q1�ŭ���D�ezJp����Z;X�f�+ϙ)�a&���$��/����wڵ*��ը�w9a/��akD��"�<�T�ފg�<� zP\�����@C+�2����7��,�����?T�apR�|�`�.�.IKO����ui^���Y��hq�V
��	�Ą�;�t�@e�i"G�����bu�	���Ӧ�����;o�����,��Rֻ5�>9OV(7�|IU�Yff)�7�N~�x��>���NS��>��]h�V�8U�	�T<�����ˑ��覮'�j2q�����|Q�������cx��P#�|�2L������n^e��5x%q��s��L,R��5�NZ��R��#YL;9�c��w��-�|�͑B� ������VWW�Sahb��� �)�����mxP�mU�3��^���9���}��ԧ�"��2�'3�6�X*J��7>
4���m�ñ���i��]��&��_��z��f�)����ѷ�F�Z��=�c�K�r!�Q�����H��� ����+�0�i�sCdβ���7��?��Yظ?WS�N��\f��B��LT}M�����n� {�����&{�3�H>�x/d\0�XS��Pd����x��'���ibkH�#��i&��H�ړ���q������c����I�lp��aB��)Bɵ6t7�<bʦ��&�@��X~��n�n^P�HI�AYD0���������#k^�.�\��e��nAQz �QP7��ѫ���������J�*��Ӿ�ZϜ�x���GAŚŋ.��|jy�fV��<���B���p�<����uM`D�p�����$�/������Q�XYY���o:5�+��73.�jǺ��^.�.:=i}ˌ+�ju�,���]mr�M���q���R��LFv�ƅ����N�|])��]�L�7�u����q)1�vU>!�Y�>pu��>R�VN�&�����yL_���$t�@�ql���q: #};�x!��~��C��ӆ7�t vLi�EB߾�K�ˆ"N��T��cIA�CV%��C��}S�GJ�Y��[��um8� ���?��dZՊ�k�����
ũ�#f�:�GGb��c@���غ��%^�St#�O���o�W�Dq�Y��25 �����:��3�0ۥ�;�n �MY�� ]70t���,��cwݘ	̋{��T�>A>+�;~�up������U_v�JO�����é��@o/]9�a�׾Q���R��\U��K�Xڤ�.�4'n���՜P�p�-��G������H�8V�٦0�(��]$p��sG�� �	�X�)^�h(u��H�v�n����%�v�����C`(J�u�ۖ���.F6|���H�ZlJbz��g�>��4��(�,+�pБ5)��ܽi^�*�����o��%��r� ��^���s�E^�.�67�u셎>Ò�����7`��4Mcʹ�0��ٝ}��O�V��M�U/�j}T���QF��l�b=�J�ҩ>���yg43U>��*������n&b���	oEJL��ͻ�b,��'%�����;oliU�I��>%[��ߗ^���T�#�Q�vO�/5&vm���}�nn*��jW���,Fm���vz���UW���@]�-|_2fs6?�wD���B.Py��U��@�n�o"��^(���|��}L|�@�h����.�*"��r�
=�ݝ���NeF���@��Z���3� �a��W���/����,ѭԭ�6��9Uq���A�QI��3�<qG������Ll9�ؖO�a���>|��=���F�mB�N�����^C,{?w��J��D�"�}�feH�}e1�D}�,Kd���?�u��,����V�,7m,z"=�T<X��I	��ۯ�]���I�\N�
��_�4��W����u�4��b�7���|X4�:1�zz,�gsO����^ �%�OH�L.��'�`%��d"�R�,��W~��Z�@��d�_� �8[>}����gw���vD�n�V�in,d�Di�w�|ih{9�5)I�p.�񽣬b�v&��?ec\�

�O�>�����I�_�����I��Og(�[L;���'u,>�s�֡��*JacU�iE����UA絘�S�.ugg�C�g��ew��?�+��J�X���um����F�U����AH��c�E9�j�=�7%�z���	��-��φT�RmY�M�����P�zߋ�e�h��˝ Psu��j�d;�6յ�_���_|�9��;�ȳ���RJt*��Y��%+�񨜤��ht��^��x���eG̦����G����5�.��))��y�;��H��ݽS`�h��p�Z���/5�����l7Xm���着1cy�)���s�:/Fv\�|�����/7wzu��=]���+��K��r�a޹4�zw
�'go�xC|O�B�h�񧼅������8������ ,�9R�����e��h�����F\�E.�[����P�8��R�Y|T������9��IL8ܻ|�O�m�.4��NF�l���o�$2���Yt�g�ʒ����7�T��fG�2V���@��?�Ƚ����v�a�=���+)咏N>�s(F�?��&TX�W�Ϸ|��倅jϗ��Wl�~��L���������st��]��&��b����qhc-�z�Ϝ���܉�I�=~���;�5��/�����x�d|\���2��
��8�H;c�\p�5�J�!@Fꜝ�J{Π�h"k�9�`bHg�q��O<{�07�]q͏e���6a|���#�#��`�Oj�,���X�Sˌ�ۀ1ؤ�e�oQ׼�"�g?�_��ju�[w7��lI"���ڡ��3.F����e�������\;����M��w��#(��2[{arѵ���أ4��'�r�z�@����bK��ԋy��6 �0����MK(���+]�{)�ol���aS�ߒ�9��G�[�g��M�>���p���0�e�ݬ޹����}��+�	\�w����6�VW�O�'��*��j��tpպ\2N��;%R�rH�:����fc���T��W�&�j�(�����X�ʼ7$��ML��GX�����(�~{���񟔃��;$;$�r�+���<E�S���at�FV��R����� #!���u$��:1@�5#�|o�����{N�яX�|�*��H�:}u2TP��$�UOVn�f�)!��oʓ��?~��eڴˣf�@:��������V�&"��[)�X�wfJ~R�;��m�4��Q�Q
�%e��N�R�:��:���������O�M�_��A���19��5x�Y�Mɾ��e�k'���nk]g`)����Bv-w��f�Õ3_�R9�^���:Һv��ݏU�E�����ųǬQUC�|��pF>,�1�d>�n��GdÅЁ��.�6��a�C>���a����^��oW� ��\O���˵TfyĊo������n�R��r�6����?���HZϩ��\i��}��ӉIl�I��@Q�������?���b��wdh�(��:�v?A~4��r�Xf*~�$RZ�C�I�?���~�<|��2���V�`㇀e��Q��rh��=���\=��Z�R��cx��<���ƈ���#G�£��m���)��Wށ�A��>� �B6vJ�g��*���c��Mv(��L�?"��i�`_��xݮ�J���8�Z���P���;b�^%�G� ĈM=�寱?(g-8쇡E�B��O���t�3�h����G�䃋3�q�Q�'�^�y�D1EC��Z;W������=C?���.>I�ϭ�n��1�a�}u1���
�Vߜ�b~��t݁�%B�5����8���Y>�*�
�-h��#�;����wz�eM�wJEC&���>��_*Y� �w5'�T҈��(�h��ǂ6�w��8q�
[[%�b�j�ݽ7s �j�8ɻ.���_Ů7`tz�!���껠aPF��|�o�軡�2���H{��E*[[V�x�B��5b�E�빀�j��*�4�[-%�ܘ6@�}�v�����f��&�e��R<�˫��*�<����X��Z\�Q�w3�ԑ��Y�Np�8�ok/�#c�ѭW޽#/v���A�x:3���(H)n�q��B�T��\_)y�f�QE����&��1��oC5�K���M�r������w���O��ݕu޿��� �ɟl��z�0�r���������l��d$�E���y)��)�1,�����`��M��s�x2
��9��[�˴���S��m�h�<���6�� u��7�v�b�(ݐ'-�$��kR��u�s~�æ�#0�)������`�8��A��&�Xn=}�/�MjY"�d���m̏<��ƪ;~D]U4qzb�	va �˧��6���0Z卻���R�浖�7�q�U��NE����yZ�|�[����%˅q�W���jB`[[C�3nf���%1��.l��)=L#�3j����X*kz!���H��Z,=0�_���O��}~�}zX�תJ�*��������v�k0�q�Ʃ�7���@����߫��dG�'�Sh�Tz��F�C:��O�~9g�=0$�!��Hx����PFD�ֵ���#���Ab_�I"Bx����VV�w��7�@wx'B�p�׳7���#77�ã�̲��}��V�0�]Wٿ6��'���`@?����8��W�B3��eQ���Fe+I���j_^:	Ǩ����lU�}�_m����.����.Ɏw�c�"㱕�~ܾ�X H��%M��K��a�=����A�&zK�i��sFb�ȷ
���T��=*(l�zMb�	����)H����**�/��M�ˍ��7��֌z����X��awԵ�ɶ�M���x(�S7�8�=���SQ���U�s��;�����T��#�u3�P'�i��	A�
q��"~���
nJ��-v��r�5���x������#�!P7�%A��]��6�[�4"��%�F��R�(׭K�(r���K�7�Y�� �e��a!�}��M̨��ˆ`�-�.�7UE׹��0_�~�{�����o�%�:�"�Z>y���y�/Gնm�9REW�̓S��'t��}�z%����{��������eB�`�曦�{d�K���4�bj���v�PRfh�a�)�_�mj�⠛iB����āWT1�%�!�\nϾ�TC���F�X:�d�y^��������F��x���Z��C�a���mOz7��H�u�ۓ��bRP�;�d��N&���LJt�'��6V�����H��55�̺�eCws���� �tћ�B�^�~��qC���P�䪎���W~��K���_%|�Jі����i$x&��fH]�ͭ6�v��ҽ�	�{�̣�Ժ��n/=Y��gM��������֛���Z��b���K�r����w�"�|Z�R4�`vu"��6p�w�ք��J;ȿ�:t䂂���qjMv��K�����`%R��ĸË�+�?�R�����Y���܈��c���@���O�ۿW�Q����Q�Н<��Z�pI��vO !�w���:>,n}����k���6Do>�AfOʪ�P�? *Q��Q1�#� *�c�v�e�^櫵t�#�5�o�����Ƀ�m���8{͢����;�	b���$q��D�-���B;}�=�mw�s&�8��ws�|�[Hw���H�T�w��@� t����@B��� ��X����^�C��YJ`�@���H�È1���cdFڧ�ZDp83!�8���H�5��i���G��v���nK�����qv)���/4��mu���w���s����v]�2[��0>U.����CC�9-܌+�ñ���5��ő��P�h�㥸��R�V��	��V5
ݑd9�����u��]������ݧ�4����z��I䷠��:,x��j�����PR��'014�e����%I�6J�)���H_�I .;jUp`(3D[S�)�}���(|˵��i����@h_��'��������L��6|I@����Y�:���ѕ���EI���(oMA��!N��i~N����:;;�UUU�,T���xMx���z7&fha�ل���a�;�7�z
��!I �L��������X��s�O�X��a��N�vSxXЋ��+?4�a����感81�v���z�ӟ
%A��ע�|m��$���:s�]{�mه��i�K�����!�n8�����eR
өT���p��Kvw���t��o�\���K5�-��8����Q�/Eha���1%d;�"���v_-�=Z�I��2mZ��,d۠�SUZ&�W��G

N���P�`�e��lف^���/g�L�8�xU<>�0��exA�Lh�Lg�����r�im��&x��P��j��ڢ�Jou�y������˗�՟zI���X���̱��`Fm@��`4����H�7����b�3�7���I(��I&{���k��K7P�*�t�B}Ek��A�۫?��2�ٖ2��sۍ��%a%<c��!n�@�/!�t�.�8�Wb�B���Ey���.�rZ�����P����"�"�(����E vm����FW��~Ht}V��_\�QZ����u_�����3�\%����蚋��Af�1"��0`�= 	��C��+�e��d���F��/DL�G7�נ]&�����ʅ����na��_y,.N���:���G���5v����_��9����ާ!ð��0���3��\�(�dt���Q�赙��2��>`���<_0�x��Y�lb�ذlg��԰�t���A�)����q��K�)&��=1^�5f�����u[f�p�θyRFB'x�����";Ǔi~wZ�-8�]��&�1?>4�-|Iu�o��΀h"��}Y-D��Y�@�-h��-+��ɩ�ƾ���?V
	�Ֆ��m���F��U7����B�þ�޿�qo����YeYu������_��vW�h�BgG�ז\0[�M�rtUU���Ӛ1=͌�FX��R(k c&\���s�vPVD�����	�|˹^�0.q6��'��kٹôz����7s,�q8�GzO5�Ça$w�08C�ݢl�7����3��J�k;�����fj�ϴ�w�����u� �J�� T���Z��	c9�2�tw��K���2��1IRW�Գ��I$��.�4^�۪_t	�T�qq��T����G����z���� �v���r>Iϸ>w&�0�\zSH�@m"��E�IӃC ^��%6���)�X��O��#Kp�v�X1'�X�
�vؒ�Yk.ȏE7�`����S���@�����A��C/h9.�BP%}@+k��հ-u4*]-�(�Y��<����B��Pci�>�2��aL���Z <-,0Փ�� 1�z�֞��0r �X�yB�:���帥>7�y���W2�f׭�ð>�q������:�4E�ei�x;6}��G�ЖU^�I;p��������J�	4�a@C��|]�e���O1��⮋8ۂN��T��T�>
35ݖ��|TD���X捲>�VG&���gRqj���#op0Z|�����B%�h�h(凤N�\���0����Q}n����כ��]��9��ox�y锄����r��	 ̤�cqF`*���b�bP_Y�UЉ�i�:����Lm"; ����a�:��+rP��j�r�\�m�x��Y
��2	7�)�5k9��`��CϗٴnG���������_�[5š���bgt�}R�"j>��{�gT?����|���7��t�z��y����;mD�=�$��S�j�i�����*�"�	5'1G�U�D�l�J�u�4$�:��"1�|W�j�d���^�F:,�8ao�#�O�8%�T���5����:m4]P��W�)�̪����5J:}���h�?�ǳ9���E�+?�q��h>q�����=�y x˲�	j8���]BYɢ������;1<$M%��6ԖQֻצ|m���8�~�R("������ȉ���Xh��l��������u�����~ ��g���Q��#Ó�v��h���29na��4�U�4�ԩ����լZ�(l�;��T���C#��#�bG��ARVl�0|�����r�c�P�Q���x_4���\�rvH��f�@b�N���ZY��Wz���KFSq/�cf��KR���W�2 iv�v��N��p�p3�0��t�w-=2���(nS_�MYu-�����h���qU�(�_�ԭ����WS����E���텵�jV
�|���Hxc���l�P_�E������z��,O��i���������I�Аe����M�3Bo�>|�Z~���I���$�wI�6�R�~�A	����>��"��n�d�[�iϋ&&��`~k���T���. XI}�����V��n������݆�������$�'��XD�H.�v��f��j=̀��~�r٦�pE��F������{<U
�s$ڛ������q�b���$BG�6�k�4�t����V���p�������cO�{?;�^le!qkPX��IIag��<�b�=:�\���o[�]���[T	���H�qD=�o_	,l�aKG�t�_C�UA�o*;���2��N�Ņ��ů������AV�v��1�UY=��1�-�#W-��v�:m��5������L���Q�!��}��p���SV#��1��
Pз=4Ԯh���6��h�`3&<Cq�Rb�ˮO���	'(ģ�׆i�������O ~�BP���<tqdh5/�"�\zy��#��0s�Q��^�.UN�p�\\:@� ws��%�go��5�L���I#��;��ۣ����6!0�G��<?k�#�؊�D#�{�P~}z~@����1YRf1}��Ń��	FwD����;��r*�<��o��=-�#��bH�ުK��ڻ����v�o�,��i�d�r ��E�����@�"�?9�]�إY,[��z0jⱐ��©�E�+��2Oj�+���q�œJ5a���dM�Q:|W�頚�����i�Fl��Z�؎�8e��i��iW�@[Oa���(h�I���UU��_ܲ?Zs�����`%��k�r���#�A��<S�y�8͕�kP�r⤿$��/g�+����h��%�[ Q�l�Z�[/������v����VVz'���ٮ7��[i����S�����60΍>1��y���/������t�V¸�9�ʾ���O��\�����W���]��o��jf��C�[�*W�"o��y:b���\����g��/��u2Yh�Zl��5𬪬̶���н��'{+|y`�A]�hcF�x�������u2���1@;'���/~E-SN	�z�L̮���@��M���F��ݳ��]�.�����p�u�ѝ!o~gU0��Ef-�{cd��>����?eɱs���|���v���=6]���؊���N�*1gd���L��\ľ�_� ������TW��G���G�i��!=|�Z),�X���{�J5111'�s��؀��X-ӵ�!�w�5��@]f_�}�L3.���?�V�b=m"�1y����㠕�֮ߺ6�qZZ6@��'E	{�MO�,:&�>�X�/Eb��9��	��Ou2,��]�j$�PQ|�t* �خb'dk��.�2n{�M��aa
��oJ���{�W!�D9B�� F��_T����OO�T>�*�ց���l�_�����~�C�����I�=�3�^�8ڔ1t�j3��f�~K�H%�?V}���RԷ��=�s��Z����e�x�W-{�'�y�wI"��Ͳ>WAl��/�]Q"�6��w�鏠[��** [�e��^ʞ~2�$��xިqf��W&��sEX]���}�C�ͣ��r�}@�@b�9:�TS�ѣ�׋|c�'�`QC�rF��O_����I7s��`~�m_W��"_v�)r���������R���YQM>�x7���ˀ��|�FGV�D�g|�~:UDe|���r�o�k�ʵ/�cQ�n��/��r�1�Nԡ����ww{���ʸ��5Z<���x7��9�!	�y��A(���3D���-ε�2;;�6C,���|�Τ����YF֑�Q�G��j���x�m���ө�h[�[��c���!�g=ݿ��T��'��&/�Z*:���b^6��%4��~y�u}Y쬓���q�]�{�
gfUo��*����oOI�.M�RH���%����wޥ˗}�_S>� �F	��*Ls=((7�(7.�&��O�����Zi�ekǔ���]�CEw�.Hԗ����*�*�O��y:��ӊ62d��L-�z����N'���f��P���Y1Ws�1a�64P���|KL��9�;؆���j���~;Q��A���|S �3fd�6l���V����a�q�gXgl��k%Q�:466r�.{q�������]����p0���Z&���d�1~d��k0Yzn$P�����+W��i�����7w7��C�ٶ��G���ͼ���BB���J�s��)�]���$*�GYn�$�pN��sI����/�ϒ7!�Q \�'yt���L��_�BUC��ݼ�	�a��o��
�؊X��[���E��ύq�������������l?��[��Hnwx����y��h�����,�v����d������Zltz��(����s�^��]&����l~�{�f���l[v�X�u�����������U��5���G�(�4����b3��Y��Bk5���	X�_!!!�%�R�B��ʆл<�߱h��6�+ϼ�{ǖ�e�i�&^�ZΏ���`~gX��&W��8r�Ǌ����]+��-�z�#E���9�$�{�(����r�D���SǏ+G��YF��Q$/��������/'M}�f� ����&�U�!��2�WVf9��&˗B�"A�&��sL��e�=��.nV�K �����?����0D咧��-���G�ע�V�����2]�����Ӟ�8A����v�2V([>���֢��-� x�X>�}	9'���|��L�Τ'�vwY�yp
��U�B����,�=T��%2V��0����ɒu��.d�v��}3�1+X�o����+������t�lI(M�n*�X_�}�>,5���F0}1z��C����߂�{8��w���U���9��V[?1X�Og�b�5͐�KK�}ﮁ{:)G�3z��I�"x�֚�Tːi�Z��5�e�ڟ��G�<��LKZ 	II�]��!��aW�g_q�};��g&	|m	��ȡ&�u���:D���o1�
_���y����ޛ�C�����Q
��e�؊�(�)�R��'��u0�˓0� ��h��}�%��ٍ%�2f�,�1��w���^����?���{溦���>�9���z���3֐x|N�,_Q���î7�.�Cb:�cmu9:�~C�X����C����C��������7Fk�"�ԷC������m���O����0M%���2�/nԌo�ώ�����}O_�0.�l��q�lcg���;܋�ɪ�Ց����2r���������gr��݁��Enc�b��,$����Z��m<��Y�p^+D��?L�j�}�/6�:�>T���e�ٲn@]���ٰ��䋣�eCw��"c�>�."|_"+q�'�4�^h2@]�>�|�1�>>��'�]���9�K��FR�Q*���Z�^��H��m��1|���쟖]R������V�{I�<�q,�Om8�
O7 4?O\ǣ�����A7o<��V�u�eo���A(���<�̾Q9�K��^��W2��y���q(3�{�J���j�i�j,vA�['�U�]?W���\�x9���fq]����τT�l�����C������p�>������5�r��D��C|�����)<2~c<fKU�s-؀Ì��}P)�TYa��m������DL#W��轿ǯ�\tgS9m�g]���^0͘���<,oH TS7���3��N��4|���t������DY�ڛ����k���m�Fnt_Qe�&y��_]͏h/@r��Ʊ�չ��^*U���t��Le�-��~�]�����'��_B �C��O������<����mì��C>�و��u��/��`�m��61�♶"�d���)��	�"l�=�i����I=�x�@�a�l�I��?d��4��D�mQ����g����j�O�F&��_��!� �[AH��s'^'���zT��AZ@*��H ���j�2�s���ǵs��bGD���.|�3J����緔���#�ܯ��G���TvX�����L<�����K�Ɠס��~�<��=w�7$vA�계پ�ȋa��6�صY�����������5��^���/�^m0.v#�Ro���$���7�L��I;�������Vӄs3ivF)4��y��ߐ�d�N��O�Kw�{�'�F�d2W��o�.1�]E�ox���Q�ŮK�!� ��[��	U�g	�Fش�e,�>�}��a���~���󆗕^��ֵ�� mbMM��^�=��S��Ʀ�V�&� /n`m��;�{���ZMc�,Ӵ��6���Ma8�2O��VʂD߷x�Dp�A�Թ�Ʊ_�O�n\��&�((��O� Ⱦ����W�&�u=4dl���JEȦ'���Zy�B�.LE��;�<��s����S�����g;��̾�?�l��tG����C��o�*D��n�ʘ�x�}|�S��ׅ�	}�2�m�*�aQ>_M}Ƣ�?vN�bY�X�E�������� s�_y�����9%�wWK�*ۯ�?��6���85Z<[-�y�`�|�{$�������:Z�S�0�r|�N`�FLKG�_ݭ�����w�J�["t���S�d�c��lZL6V�T��B�;��0E�p���K�׆�_����=UUU�d�io�d��ֳ��^	��ӄ���ו�ѿ����c�g���S�Qh���̋C����ó�x���|�h-?Hi"�����s���K:[��#�M��V�CF�/QXG�k�J���a���"��[&9U��w���w����$'��A$]߿�^�u����)y/���U7�yی����@ANaa�~�����ft+l#�'D���kX�����f.r��>�r���e^Q�W�╒"���-�p��i-�E浡��s�!+����G�<���K�7T�ϜP:�����V�nK$e��昘��n{D�	�B�����!�ຉ�5�m� h�m���#A	���Dl �x��A>�N ���f�H��T'R?]����Wo�LsMp�T-���� O�|�Ge���Ӷһo����S��C��Q�m��_�Ը���G��r&��B�@��Z�A�/��މ2��Y��ވ�0�!]Bғ��i����gnfx}�K�K�y�����c��K�hm
�A�n���L+/Do<d))�֑��j��@@@�)�.������?�m��c�z����ӭ���~�[Ì`�ba0��i�"Y�k^�X[�K�g��WiK�1���	���foД�.�+w�߶��~֛�jS������.�Y�5����)�s���G�4��%B�
�wP�=��[�^� ֞�ޭP��T�]~_j��Q���=� M?�3��I�p�f��z�D?WGG��n��k:D�J��Ҝ;�7	�����1� e�l�q�Ug�:����@��N�#_�|���v�'N��aI��ܖ��.��8������Z؋B`�_X!��rˆB6T��=��U��˕����Xmʼ[�}sޜe��i�`L�
�W#d���k1��p��L%s<ϼ]�O�贋]����!��8��F~_Y��Ʈ��p~�c�O�<���o#����5��]������� /���T���0wh'h���dg��88:;+�|S�l!j�9����û��Y�o��y�=�OvW� W�����J��[s7
��m�_�9��O�'ॅ/[�ȼ�?
%�#����Z�`ԋ<�ɩ R4tAa!Q�f���V�-���3sss�t/�ݽ{���c�`�5Z��-/^����O�D���(�B&DU_Br|���Ĥ��!{{�����T��A���ۓ��ߚf2iV�7��c�S5ս���[G	Z��No��c���U�5K��x��̵y�:�c�п�`?W���x=�8���O��022z�1�UV&a���V㎙ߘ�����������R�e7�"��LO�3����ƀ��}�{5�}�H����ɕ���� �T��@�Ļ��ޗP��{���"���je�|����6�A�`,Ex�5�G5�vU��}��d0R��Ѩ�ܲ���3��@�j��	�,*��os�ց\��g��6����b��q*��
q�����rS3#�X2��b\l<�oȪ����B��gY���!;;���Ot��z�����-��-n�����5S-�-E9��[ה�5��ޭ�q
�����2�ESM���5:�������(�_����Y�2��Q��y�Th��)O��m�I��G���]$ΗUP�(Y�ʊ/��ߪir[�D�v��+W2�����d���V1�R�=�����o�R�ѐ�uB���*��O=�Mj_YYYjhhpأ�)�9��z*���.Q5�H7�N҉0��=��z�@{��|�_GIWg����\[��i���O*�	�����#	=2K���|��_�1[P(e_P����===�7n�0��/+--U�;I�"�(�ɹ��:�J��'(�ɰ �������=�0�0���;�k!3��T?�	
�E�t�o�ꘖ����U~ihh�[�1y����WU��26�G^^�����7����Ú!����WϳcXD���.Xn�Āj��������,#痼��-�"F,�0K{�o�q=���-�g}�S������wK*z�\���s�X���d�X��o�YN\/��&>�eiB���(^��Ǐ+�����l��xcS�����---!Hȱ˯��i�ئ?D���<���d�1��_��ZZy,�����	��6'aϗ��mA2�[i�'Ξ�_[WW��g(�F�IKK/����,� <���V�G�K u�9v��bcc)�jK�#�m@���Q_7��! kj�M�����u*��N���&s;;��W�Z��~�Ctf�w������3�lқ����e�?���=�ؒa��2��~�PU=z�hUC�g��/ �l�O_�V=����Ǘ@���dCd���$�B�|6�,��n�~~~���l�GS��O�QZ����������SIQ���������l9�V�5�I�k�y�⮣����EǓR��X����'�O�w�6���35_"�����%�|÷��i{�x�ڦ���
���ʩ���F$:�/����h4�:f�B�Q��O��m#k��噧�gyޔ�Sަ�'�I%+R��UUTL^�z�u����~~�Ϝ�i�ܷ�\��'|�^V�y�4��cb|���DE��3G�:킬r�f��14|]�:Z��D�"�K�|YqP7>>�~�e���]%{����n��=�h؄�/?�Ϸ_Aw�<��&C4�j�UL̸)	i���c�{{{O()I9`+���m�I7�t}Q�t���6��i�e�t�sV2ژ��$�I5�g��i\�U�������"������d�	���ݴ��/D��Ox1��?�D�D�9����|���b4�|����֚s�j�|C:�C777G���	�3FIRC��֮�{99�|��5��@�FI.�\�d?�'����ǋ-�A_���E�5SGό7�M閌���M�����B���uit=��[�N����,����D�aX\�}�������03^�U4����}�mC���:�O�]=��Y�cs�@���6�檶����h0���!��]jhܻ�Y4�W0[���[]�J������u�|���@=�%����7����>K@���݆���舰0��&h���U�D
ZXX0���2�/��Yf�d0��2��V! �����
b/���,��o���y�i��d_H��G�؂�L�+ϵ����қ̻D<v��̲�+��Nm����U��I��k�<��~_+M�jpS>��Rt��I�Q��v��O&�ԁ�E{ ,X��pE�Pp�֑�d픹LP�s/r����]�.�W#"�,2C��9��5�09���yݵ����=���$Yw�2� �[k.G���RY���v�"����>2��k�K;R�#�3P:��Aà�1"vmi��k``�ṋ���?�	x�;��\�c��iii�=jK�b}P���L��X,E�V��K:B�΃~�
2�E�V�֬�>|���K�6w�����!s�C�O�'�ye>�{,�䘢q�}^���+������2��:
��zZg�{)�&�;w�xS��L�)���~���0̺Ѹ�pB���O7�$VHZ�]���{$$���i�Q��ϟ�X����o��5�jv~��~u��2��$s���e�/ӝ�ɟ�����gnE�N((���oBd����z��Ӯ-���Q�Y��ȟ0l���]��ֲ,�up���v�g�Tb�J�ɪ.|�1V\\|��܎���Wh&�������o9�`u�'�5Y`<x�r�Hdz�}���-j����}\���u��̍��0�E��b����Lװ�A��m� �,1��:B7�����W]�J�
�LMM� hٞ��?���#+�/W���~��*Id�9�g�'oz�^�d�FG�P[$c�������g�7�	K#c`��dj�-�*���ׯ}�rrN�Uo����8�<\�a��eB�)�ˤ�Q5��ϟ?�綨
��T�v������l�j�K|}���,s���4��7~��Z ��$�"4��`/"���OX5�L���m=řB@F)&a�#�����_�eKd��q!��78��_�~�C��a������\��4�@X;�z�o_�B'*B��b�ӹ���k��X�+��uA����"���aQ����
�g��м�1(��~��)l��j���k`�:	���,���܆H��S;�e��5�'Wfʖ)�=�[��&64?�"s��H�pF��5f����?[�kQ��zǈˊ��Aa�x��:,ܿ�od�z��>:�~ߕ���3���%�o���/S�[JPSo��f�T(�"`r�)��!�1���x�x�t��;i�����J3�Y*?4�ч���%�2
�օ#yY�Q�c�эc�N��=�)�Z[[3�IW�]]��""���J�i�Aa�̻������`{���re^�E�k���K�y�#�Q����l�?
��DL/KD&��x��z�6��7��R/- �����?8pY8TGқ|�0("1�GK��A����q��cǎq��}A�~�?�*P��e�Y�P��y�:=���mn'����b�G���x�@��6&e}�;�D�P���؈�oT,P6�����JJ|�
��;0?�C���ߐq���AO�@�aFҕ�Q���E��N2��vV�?��<��~��^����PB�*����2O�fR�!�AԐ�k" >�P�j�;ٽ&�]��z�#��C�]�2��Ξ��v�W!��.���,ң�4�y��<S��{R��݅���O�OF��h�c$�����	�:)��Tr�|��J�<[~T\\Q�<eU�-?n����OEJqQn���ԛ^�M?�?&��Ă�K� �k_]���#[rX4�\vb��Z�{��G|��T�&�[�1GW0�4�4�Ӈэ%6@��j/_����p��H�)*Z� V�X�G�b�G�/d�29�L�}����.��t:�Z:ZKPD�*���{�S)�����jgJ��ǓX,n������Bܬ'�
M;������V���̋jS��!Ð睖��"(�w�������'?��c�k��Ø�
"S34:��r����HP͛<�Z[�![��
��k���$!sRL�MH��	@�1�xV����7����Y��o�W�h��^��~�?f$7�����;�XzՐ��Ffu)�P$�x(�gP����p��sPP���#��1�*8w61�nJE�񫕙�ʼ�
F΄���_���ƭ��x�ǣkW�����0x�:,�r�ɓ��!�J!e'�wz kB.�H�08PG n�7�	z+!�=Ю��S��m���n}[�0����P�T�>��ccc�O����	��D��{�1h��*<�C��خ��,�!�,=�m��>j�N��n����>��'�dq4�9/��5�3�cno/]�f��555����:��Ӗ�<�l�*2d�-\F;�f��Ud�I~�������!î�☊��C��4Q�B{�b�2=$�L�z.S��w &r_�u���& 9�H,����Ki"�(C��X+�=Y�4x�|���m�x�"�ԛ�w���������/���t��	����Y�aQg��+�Uo��Xi��y�`\y�;6�۫�#D@�;��d)	!K���UTD� �� b9�����t���x�n��
����q�r�
�C[; gg'�I����}����h/��]%�hݍSp:"�k7Ax�B~��F#�!tH-����I�Վ���\�Б��>�@d"�����S��{x<��bPSd�ʅ���H�>�wޛ3�Y7c���K�����[����0#OVv����u��aF�0����$n;�fn��B��֨Px��7��cz�G��LKs�>�1X�t��R�.:������]�	�C�(H��!��@��"K�K<i��MJM@T�;��/+ڈY?�qh�qq�r�[,�!����B��/��Z��+��Ϸ�K������kF�����Gx����%}��Hd&z�����Ja@ѩn��B��Qp���rQ¯�į2���״���ա<���Х=�#*99��j�u�S�j�x�q�߲��B���E��߂z��M����U�:#<d*s����qרm�د���}8F�������l�9�YU�{�nF}�e�q��(����4�1ײ�w�9�N$�Y�'ȢP֚	LˈC˦����@� ���M���B��WM�2��o��-X�Xի�wQDERJ��mI�*�G�W�g�G&k��4�{omL�؉��&C�kd��^��w��I$�P�%���>���%�|�?3����ÿo����7U3"��;��O525�sg��)=V��Dk�a�
X@X<�Z;�}�_��e�v��m��<�}����^�x�xB���ޠ$��Ŷ�յ��	�3�~B���v�F��m�hm6��W-���q�����\ f=��3�oH%��u.:����$1�`;��pdj�c�Y��u����r
)��H.��ֿ3Dn:`�!۪�`Pg��W�hF��p�6VnImV(��"�#G�)�d���}�B�!���`��5W��֮ҍ(����A�_y���G0	��;��r�g��2�|gYggY�l��Z$ȑB	g�:
%�-Ϭ�25!H�W�/�2����hg��$B�H�X针���ځ��j�*���.F@�g� �׌'�*C�Q������N����~�O�L��Ner���GN�y�r�.�o�R���CEJ���8��H]�}�+���켺��ā��Ql�z�g&��}m����͚�8H�&�=J�^b��^�U./D�z�ݜF$����Y]�}q���d�lgd�3�5գ��J�g�����Y��{_7Y��7�Q�8�����2&%��m�����:=�)�xѳ�����`��e<��b�����Ptj��M�B��"�Q]��_�^��mb��>�| \��s�c��L3��3<�.W!?�ʃ�RNN�&ܐ-��]�{{{G��<����X����$A��$PHC���~�Y`ݾH���冇���`AA�4�{�I�~7�����98:::E)^;c�w���j��R��W^d��~�Bd�mJ�Ą��ׯ�EFFF#�@ï�ῐ���ɭ�=�Pq8o�$�1X���Խ)�ʀA]�1l�;���[J�sCE�p"1�ɓ'�3�ip����������n�|��n
Ad�!Qo�����1++�i�W!BCb�Ԉlh?S �����{�;0 |��67�����O�>�W*Z�m�f�%�iy7�Dy���S�W�Dܵ��V��� �|?�����W\87��	��T������S<�P�2?���=�EF�����a�b;��x��}������ �|�%2G������!���2��j+��@�!�א�gdZ��q�>�~���tҧb���jO�@7�xmk V�;D�;���(^��������шv�SoJA����n��&H�|�v�F&����|�<�˼L��p�Fǣ
^X�l�[��oɮ�13s0�;�'����w���z�@8(���v���o$B5��U�畔(M�KE�qG��)�Lµ:(T?��{��K��!f������^�@��j������p��0������j$#��/�ݖ_a+�"vQ�&��N�4Ϲ�n��9u ���{WQ5Ww7(>�8�����'h~�O�-ms��a~U���r�y��,�����q(=3��������t×�O���V禋qg���(A���F��f�R����d��)�F뤇`N��
v��8���!���e:<8�ś@ �8\�'$�@y�#�&i���<���P�\a�q�9D�z�{~�e�0x��N���~~�w���3q�jQ/���YD��k���?I���/�������eW��W©2����"&�*D��}G�#7꼾3}��_T�b,���K@��i�����w��f���nϻ=����=��!��'���Պ��Fx/̄l��W҇=j�*�ݝ��&�)���������!��>n���&a���s��*�U���U������ͧ2��ÓJ�>��7R �,7��:rQw��{������ u]Ha!�P�M��]�3�����fˠ�eo�ބx�`��p�@��;�$D��K�b*.��	�N�er}��.C�R�	�W��y�*��R������p��$�X��8�@	k�n~���Q��*��糩�{��o*01�:�k$š&�J��e�t��Y��KF��sk��k�;��8��FT�1U¦�}Z���U���2�n�dܣi�U�c[Ά�9R�䝕��S�E���3�6
\y���c$\O�c�K��w��}~�?�nR��KO�kPOI���|�P�� �߯^�U��"���nk�H�OvI��~g���,c�u/���<��c}ff.$�{/�>R>�h������w+�����W�u�����Y�O��W�_���W���s>=-K"��7-j����)��%�G]wQ)�!���z���ס�M�0��ò]����V�p=�J����/YH]��F&�k%��ws3f6D!���I�P�ݣ_T-��fd��d՛���"�\�:��s�������k�����ɇI�'�pȽ��555�%B�9(8J#��MV�NN��/N����A�[R�����5����H�<1��y��3�i�wk
~_��盜��#��wf;��qsss~xxxVv����*-���#=Z�Gx�#�4<��5r�8�B7w� �ٌ�y.Vl�=�.aw� �a3��IK����W�F[��D$q��F3�a,��4m0|��vܙ�҂�}]��hd��́�$�_�6���?�>��215e�'vjj��9��!s��i� ��EeAnF�f|||��N2�.�m�gdY�EPy�A��g\�{z�N����6d��S�h�c �c �d�������٥�vuC�����+���188RY&�S���G�<faa�[G�Ef�9��[oo�n��m�j�$�������� ��w���ʘ�SB&[ǼxQ�+�=�4������ǃz��/����vw+����y��E�(�����������14�%�����ׯ�����)����!d0t���lȯw���Ϣ�`d�&&&��ň�����q ���=�-C���ff:ۙ���Q:��Jطo_������H�a�[���ǑO�>�uum+8	��ٞ:`��_VV`�ƍHs���dO���rM��?�h��*���%d��� sb�&J�OXL�q���`lb"��\���<bq����
w����qJ�v�lmS�b����Q�-�����,^!$8��i	L�u�����A����bd9��Y[[{b��w/z&��Hю?@X' ;��u�T~������+܀l�8u�)X��Z�
�=��%���67;�t#��k��e�]X�˞���50rv����::!�^������J�\��8'TTD��>6Bd�j��e��O.(�O��766Z��|�W�===w0�SQ��*DgoJE߻{������U���{#�ի���+��0�h��H"�#E�(s���p�),z��g	ɖ/%!m"���oz��m[}}��ӧo-�A��W8}z/�8�F��'����ü��T�}=\]��0�߆�[�O�EH�wLL2U�W�{��a��s�8#+����>Y*��ܫ��x5�WC�N�R�Iӯވp3�տ��ָ}�v7��qz��_Uw}�z�%RHHHZ����#LF��"�%�W�l�}��cC���m�?b�ԁ�|a�Y��!r�^���:_�㪌�o��r�Y\&8:0?��2.��?n�F�Q �蕔��sqqY7$�G��p=�߄3������1�W���ս{^�v-hll�@�mck+	
	IMM�>P�=�O0I־rI2�I���b���xp���#q��Y���l��1��5�L,͎�Y�D�����e���^���8�Q�������͗�_K����z(I޺9셊��$):��wg���n�q3�f�mS�1������2|���Z�EE���?�8� ����vT��Q�^Y���ԛ}��{8V�#ŝ��1����k-�_��������C�	}���OՁ�`	(5�۝�$�Uts<��fs�R6;;���"^F���k�YN�$��c�
l�y�F�gv�n��e[�d��MV�����☦/d��3�~�Y1��[2;��I��(�{�X��=5���a�'�:�_���r_�@13<"":���c�6�,k��D�0 ���x�)X�o�<=�0�+sz��M���t���N�����x���<#zk���	����Xb������BD!oْg���
����j��+�Z���_�QDr�chD��)h'K�@�����x�X����^p���{as��y%�_,��u/L��<i���0���Z@Q^^^���L�D�(w��u��C�H;;;kZ��C����zd�[z�,�8�dCK� Y�u* ���?��Ssp8��ۋq)DC�w�$�~�È��~��P��w����O��*�oc;���X�j.�]F�B�zm#�Nf]����s���3	A9��������Oߣ�6���?���9p��-�YD�"""�z;���R#c1f2�c�ʟ@|�"jB�z�Rˌ�r!y��+C�%%�X���7@�  �ԓ֥�YPZlS��R�$d�8�B&è0tn�%��-s}(����8H^hM�*v5Z���a�8�h����Xŧ Ԟ����N�ⶢP>���׼(:�`q��$��z���4�	���t��g��gz���gy�[[[o���9�.�V׽��52ݛ�V�Uy;�%Lt���<�e/�.ύc��9�Q*(��Ф�d��~���-�>vN����ݓ����9��;m���w���b5Xea�߽��&:��(�|C�)���kI�,,F$���0
�1��9���@ �M�/���:Q�!
 ��%��U�''��N���˜>{��o�+�'Ɇ* �����y��(Ld���(˫�4��ب����,���6�5�?P���Rt
�Uth�-[�Kq�i���,��Z�'���x�yj���ӾXh8p�׾�SQuE�7
"d�z�^���p��BVy����X�5F�Eݔe˭���xT�e���wQ����H[Tj��	�{�K����Vll,��|��Sژ�u�����V����OcB�����zl�Q|Q��!��&�N�ܐ@�*W;�imf��vG��R�ߍ�f��Қ`0d�ȹ�w��ʆ {f��8T4#,����3]lx^����b�ؐ��+�*�����߰Y�eK�Tpp�{S�`&^�:gL!�\����AV����3�~de��|ͽ��F��
z��r6)���G�	K�^�$�ʭ��&�����2��Db �/�>���$a`�#���$"8?���@mmm�&�����
Nu}��,Ҧ������)"���&&��v��W��X���x,D�R�c �yy-.�������H�@��U:/EТ�г'�+෥�1���Y�v���T%`m��^Y�	�LE�߿L�P�Gɰ�� Ml��N��	������u�[M�Г��B�A �.��|yUl�ȋn����ʷ���Y4r.[���H����s��~QGν0���{��yIР2�`���&����� ge�k�+�m�;k�{	�&d���)�u��.��@��{s�!C�m�.
ϜI�v��a��&r�m,%IgTT����~�C�a�����z�c�k�8���ʡڥ��F��~OrY˨S?}���|�$���3D�Wa��q��$�̭�c����Z�
�c�D�7�y��RG-�0�}�#G��w�f �!]��R)3U<����$W�B�D������9�겫��Y�b�����ﳸ
T�;�28X��/Baz3�|(�Vd��bn@r�� ����0�X����2�y۬�V�>�N�]�*X��1U�k�mKD�0˖�)=3F����� ��(������2%��*`,�j����]�r���꧹Pk�Ņ���"���D!�￮~��\o�	yВT��k�,âՖ�F�R�i��x���AGG�$};����݃q�>'!'�R��xË�Q�$����m Fu��nd�+|���n��ZL���F9_>1Z��o��O���*w�Yp������<��\�A`xJ8ZW��	P����o)����!C��p������s�I$�	Hv���2>~G���#����%"��}θ��

��i��˫-1���:�cFO\���`Q>�f�-�XuÃCCh ��qj��EF#���ވ wG컪J�)��QZ_��h�5ȿv˖-Vq���E\����oL�����Z��=�_��c}6�^��������/�5Mf�iI.̳X!@��a��T�����3^_S��Խ�|3�o�(dȉ�`�[!i⻝;��x�O\_g�b��M���f�O�ݕ]͌�0J�q��jecT4���bc���#$��ގ�~��4VT;���)-�q�ҡ�m8�:rTG�T�陙!���Y����>C�I�$��p�T������(w�eI������� �d�]�[?�Q(�ʦ�����d|1|��r)�$C�����N$�AZf��� /�D��LNn��ȕ���H����B�1���h�MC|��.��A��uO�0\)�����\k���C��|9T0�2��37�YT��Ū�_�d ��C�{��MVs�����SS�LLL��X ��3�/d��tڝ����o��wD�^�(Q<��}��������T��n4.Q<�~@��Q�
c�^�����/]�3:_�?Z#xAw����7@O\ ����iF�녳EllsGz�A\h��{����,�ﹲ�խ�9��]]]U�� 3wT�Kj8�XG��ۭ7�}r�^�*�J��H?s�7ڙ0��\W	�q��Vo��-))�+��Qf7$���Axh`@�t�z���PI�\�]��՘YR��9�j�i'&P�����8��۠�?����}z�%�z�g=�~Yc�[N���A+ذ����=�F�0׋XC�"��S�/˵����?"q]��4ʻuN��g��YƬ��g��$��N�Xi�wzژ��,��/IO2aF����Ƿ�����e�^��1z�����m�J�M������M��&�w��(�7]�@x�t�^{��P�����zZ����>�</���ZG��=GlD
��3t�l|7ۙg�U���yĮfc�d��3،RG�"���glQS�.����S]Wٍ���of�O|�>�6���ٷ6[08 :bl8_���$����)�/N���n�IO�
��Y����5Uǅ�ͭ���l��Pg���؞�ʛ ��*ߐ:=1уL���j�zf��Y}��l~����p�¿�c=r<my8&r���G}�TtC�:{�����R�!���:�3��f0h���B�`��>�^�&��(&0�������\���BܖUGV�JQ����J��hH�)ooU�~렡�nы4.��B�����A�Ҍ~���M'D/N�+�i�h�ڮ:�/%��*2�1"����3h�e��2�o����\��W�/Z����u���FY�^�>I�zLT�!\�ϳ�a��[Ϛ>;l���b��5�ԚL�R��D��Ñ������E��`Vvam7�����X����>�����n��g�����KJ�2���_���hH�쭄Ѯ-q�4����n�-���tf��&e��������%B)F��(�p�ëPǨ�"���1�>o�G��A�ti�<�!�gï�-I�!p�)��7��2�T�T�{�yzd�V��pv<�ҷ�j�E~˿���=�6*�]�B8���;B��'>�nU���zO.)Y#�V�}���Ca�g<>u���M`"�
RF֔١O����*������N��9��G���vT��TV^eK�֋��>hY<%=���^���
� �|\����n�)���n_�v�~��BT;`�o�(��1�� <,lի��9�G��_c��gH�П?���~��4.�+�t�,�xq/��5�SSX�]tq>���|�mU�1+_��X|
�����p�1z+ڽ�(����̓e�! ��zZ�n��� ߄�[�S�p}}�Δ�޶�١`~B�*b�+<�g�l~a���ë�(�i1&{��+�q�\7m���N�����-P[rc3����!>w��.��A�[�4���7�,��r J�Ҙ�Q�E����r���DN�K�V�s`�%�`���B�#�I�=�ɴ���6��)��ar�6V���D��_J\�����X���$"�kh8`9��u���(RVUY��D����5��@/���4?��l'e*�6�+f�\<��_2P:D#�rZ454>{E��?Dk4[�����ky�	ySrZ'��u�ߟU{�������ӫ��E�X�i8�-�|2$ ��Qpӑ��ե�ެ�oTux�P��Yf��O���zr-[6Z������&��8�n��4�ڄ�G^@0^��{bP��.��0�.j߽� 6�mH��f�~Q��C��`w[����#�V�q���j�P(e�A!@�!D�`���P{C�DY�`i�Ul�X��v��yLrG�k*���F�Q,0�8MN��Z�+W{\��� ��<���ek��%H�F��סK1�BЖA��/_�����!�PY��ڽ�٠�	{�X}ߕ0�c�3HB��x��!�%D\PTtm\DD$@,p���e�<�D��Pw���@%B�^\�^���J>@�!D<�Jdq�{������6��B�P��Wv�)���ͯ��9���{p!S����ё�^E����\L���?F�e�����#<��;+�YHN l($W�.^��#c�Z/x�!P�{r���^�%��=���'FO���0˖�!�{��kw���6����*;���EP��5IR4�"П�H�b#�������f�����ոͶ���9f�Se{�w����f�!+�:��(sU������[���-�Ф"A���@�#�-Ȭd��H�$��G�^�F�澂���&vi���ͩ�_A�K�^>�LE�r�,��#�C�Q0�B�˘~�Fd�,Q�4#�s��ءiS�5�� i>R�v-g|c�d%a>��dk��8���
f�t��&��3����=�d�J/�7S)�T\�j�&��Vui��2w��z���U��=�b�X-I
h���n_WE宁�*K�q��+�x����$=�C�3��#�Q�A��<��[٩`B!3\f��U�>���ڈ:':i�.nV���P�����x����B����>Sѕ��|�c�bԸS�&���[$Ei���Ъ���E��@�"yD���Ń��:C��t��l��,�q��}�3�@?��5�ո�u?k�~�d�,2��%�����ǿ��8>���|��;�^��~j��`���	��_��&���0�kid�$�1�$G�⻵3Y���:J�hG�>o?x��ꍕC�VKX�Ͼmp<�ʏ�W��E���:tۊ�8^�����a}��]��]��/�j8��/�8�t<�O��p�.���:����=-3��6��'������[t��~���ϩ|�T�響�'�f���r׏��t�^���)�3�	lw���\̈́Ḓ�TwmZ1F;~n�>a�L�0џ�9�-��-�}J
eJ��א��Ul�l1�Q����.�z���n,nn��`r�>��J/6�W�	!:!�/����$ٱ8⏸+k�ǾSF��fJ?�E�������Fm���Ct�;Q�6�����8��]V�a�?�%�+��࿂�
�+���I�]��s-��(6�~����R�W�S4]%I�x�N{{�ݻ*�v�(� �2���z�N�ۈB����u�3Ǝy��X\��皢˗�"�aKY|���V�<�cIR���~;&
�%֨��$E���oܘVf���lG�8;������ʻv���/��Vꜧ����[��������wh���!��ό>��xH�}g��>h�`>���4S��%��.F�[h�H�R�#�5Q(nh��_���K��Ei)3P4���?&?���Xb�'�����5��z���E�|�{[�8�n�MU�ڻ�@(Ӷ�t�[ag��v�-YbEΌj4mBQȱeC�Ð�`Ȗ��N�uVҬcBcJ�fDN#3�CLcg�w?޾������������u_���]���<❳�����*PڕjW4ڠ�! xy��=���L��^ ��H�"�s[ ﭯ� �{F��W^l3�_�y�b̅���F|�|��㣉i������ѷ�I�m��t�G;��(�Nn�Ȇ�HA����~?'���yʈ�	�	6E��F:���������B�
�R�e��#;�ޙF�餞/�ZO&�,�d�c�l�$��$h�ѡA�s�a[ K�-P"*������XN\sW��[�SȈ���n�ڎ�R��	\��QjM�������Hԛ�nB#�u')�F,�ð��@:M9&DO����ф�a�����}P�O�8�[G\�D4�q��a�O{ o|�����u��:266r�>B�$>�PB�(���fBգ_�VV��,F�?�7��b8F��jvOV���@�>�HҪ�1�8x!�鼺	��C�/"X,��E�R�@ ��*�o���Gϸ�pis��tR}��ꨬ۝(a�J��葉��g��������=��:|�p��&�m�#�Xcg�TdA9�  �!(�tC����S��Aˋ��?������Q��?Y�Dj����q7�� /t@)���>e�r���&j��^*�݇=Ã�x��m�i��+4������HD�y��SE���-Ы�X�Np���f�����?Ny�x[�A����-	^�MbSz����-g��7C�-�	3�����B#��? q�7��a^Ƕ;~��b}^fVV�O(d)#�;v[ʛ�� �d(�"�>��	�(Ѥ�C P!]��F�����@��fO&G��Y�	��q�m��a�qcc��Ag�0A�AI�Q���t׃ϟ9X[ZY%u#_�;G�<@�xqX��pH�/|h��5�����)�W�����s�U��,�}X�[Ee��Dr<�E���-hq���F����Wo/ۋ�k��<l�ԃ̬au��2��	�H�҅������@^��J<�Bmj0*-l��JR�6�Dv��6�0ݙ�4	7F}h��66��t�*1'�X{d%�+��N�60մ��.��!H�$8W���Ʈ�[�w��:o���s�w	��+�K���1��������D�fk�5�+q������'���D)��_#/9����%0؏���-}��He�@�w�s��l��&gQ�z��YM�ò ��V,��Q���F����:�dV
[7��Yp�M?\<N�� tO%�cA��ޜz�o������@�W�]S&�]H�|�WfCP�4��9W�n'~gw0�a_hP +@���N|�Cxt"��v0�� ��Tp�@��qZ��7�>>>ƨڋD�֑�p(O�2;�_�=��x�E9��k;��#:fi9���6�	��_����A �B���KgO�
s�\��Am�a���"�U@�n�M���Z���׬D=��n��#�Rr���9%�å&�ռ�@p�Z	���?�1wqq��ى ANH����;�B���	O���v�:=o�����
�P�ݗ3\[��E@����ۃ{���S7�VUUe#�܈Rs�YB$p�bFlCzFF�aA0I��S�2=������ڿؼ�q~&yLR5Y���=W��5�H�u>�B�᯽�u`^�����Y�(0�՛���&�2�@*q�9�	��c�F$q����Q6]u��]��;n�]*l;k#�Ȼ���2�w&H+�m����SaF�+����V���|B�<{���Gg�1�F٬$���%��8�M�S�s#;37W����7���� d�Nѫ��N�488�M�tT��f��|�x����;j�'��|ݘ��v,���_�Y2김����|�����rn����P�<���3!'��E�E���Q�
Z�#�r���H,B
FUcJ0���Vm�f4�b7�g
�ր>Ʒ��3UJꄏH:� [x7�/�E��u<F3<+�7�I�o���_�S=�p��#�u�Fz����dh�NPB|(4����xg,�2�,�T5s6AkXX��%.5c6g��{������!<��L��T�}dA�Y�1�S�c����⮶�aK���E�(	ň�5F��N�Y�.,�~bW4G:~��:��K(q.��u�K&#6.go�a�*ņOs,�M5�	�}k��e�H�h=}ii$�Y��~K�X����L%K��R���a��(����|v|}�#�����3���@�U�*�]�9�{��M�K�#��Χz�5'��)���\ۛ��4T�-�K�{K^�[�F�&�fTl��x�uS�
�c�C-57T�z}r���S�(��{WO�	�@���]3���M���n9��R�lR��������LX�ag~��jF�O��В�/�	J�L��V[9�IHb��l��uP�@�%''���qAg��+�<6A�D�4̴GSf��پ%���e�V��ߓ_G���}Wd�dE��ߏ�bn���]&��vZ�E�_����x��6ы ��$	��WU6C�oA��ac���_�*�4u+I�i'̱��NU*�L�}���5zV����\��#�i0������,��D��ϥ�� TGoO1Mq�V�����2ui8]�0���~DY�x��=b�'������ܨ�r6�Ի|t�_#�me�V�J��-��*��ĊV�O|�Jy3�f���&�k�Ô�^!������i�����,:%'N1VQ��Sc7A%�8��-^�S�R���v%�5��Hٟݺ��D��݄�n2��,],���p��2����c���m�Ay��s��BԍV�$yj�����Kfш�+��ґ��o���V)�r/75?I��xt0�G(_n��M��hT�WxyE]+��Jhv�����
]��뉓����F{�]gY��Ϋ_?.�1�NJ��M�mm�-WL)/�@۹1��)Cc�y��������w�X���ŏWD�m��O� C^�/�~@)a�P�K����c��Pp`8���%PB �J��e�'�X���C���v�l#d=b�ׂ?T� ����,P��\�m� Ü?� V����sX�!����ȺW!HV�. �`��k���u"E�i�=�*6:>��Wy����M���_tTԫ�԰����F��,���{&pi�L(9���� �4�Jb&�n�p<�����hG�A%uq7A?y�8�y�8��V�~�D� �|���2����+�`���'!�ZƼ�	�Š^��HS��L=el
?��/j��%�&�&��T�/���;�)7��'{|B��?���y���,m��`Xlu�#b�zb���[��B_�:�[�>_�Qd�M���_s���zZ�������|T���v�:/�h�������o���R"���ݑ�k`�Z�U�?�� UD%%�do��4���#����r|L��J����-�M�.��=����gs��2��Y�Ϫ��E��4��ˏ��t%E�2����i�����U���)Q%r7ݽ/�"����6AVp��_N�@v�r/�̼l����lLѽ��}���Ge�8G[p%��j�����n����<��|$����h�L��MSjі�e�H*a�5�,���t`ܴ� Vv�.��s�X��r�y9u�׏*P�w(/1n��~Z3�t\j�������O�&�8-1�>T{i=�x���Ɯ��C;�Is;�n��3-'�D���!#���Bm���Hb��G����ty	B��}̪Շ�qM��ziެ�b���d���ው��zf�և_�؅O`��j�.�{���_~�b��0Q��Z���<�F�
o�����[6;�2�w6� 6�����M,�6�6�Nq�K.ڙf5�E:��\��k�3˪�{��I�PQ��j�T�k��cͧ�~��)�ȿW�A�w����I��mT09B��v�`x�E��
�X�?�V�9�{�}���H��rz�r6����OM�����u�,����n(Oo��\5�����T��T��D8T!y(N�0T}@Ҡ���U�5��z�Z���
I\��p*�:@t���$�4V��0}��D���r^If��j���� 9d����m�/	djM�x(�(�����"�e>"�T�Cw��~���WZ�����l"ȶ�9�����K�>�XYʢ����;�]Q�v��1f29d�����3R2\�ZsM��>�Oa�?\b�@���17g�B���7�����l�DCi}�uS����Zyo=�q,DMb����YY��D�b�(�<�-M&���8��"pg�d�o�cF�~�n�B���cR0���N�(By��?&<d�w�P�,?���/��V?w�-�\��TO���C�&�T}���?'��)@A���)����|n�'=�Y��P��t��h�K����n�vh\�;�]*�壇l�1����Qc����bȍ�ڬ�D�9���
)�}1�o��j����K�K��E7@��2Y���� e�1��]JFQ^ؗ�-ʹ���7��f΀z��;j��ϻ6��-��^\@ˮr����� ��|�p�Ej�dM�iV���0��U#W�}sFe���qٿd$���WK�f�r�e#�n�������
�����3��Y���'.��Kݚ�C���G[�%�4kyx�5�G"'�6�A�~)=�z��ο'��B���W �? t�e!x��/Z(Y*
Z��N2Wl�F�7����z�S�����ݛ��0��3^,��;mEb��p��b��2��춤�߃Y�y�g�9)���i��vt4ׁշ~���k�`�e����� ���"�!�ԕk�AZ�<�.zu��}�M�k�h˓�a���kK�Dj�"}u�P2S���jO�"�P�^�&��;.x�!y�ݏ�T�!p�R�+���*l�nX]s	�)>��K�T��U*;�L֡,�8Q�Xg��v��w��
���e3���;ү���80uPn��{hP�N�ݽ�.�s��<�s�1��ڃX��[����l�]�(����\�#�l�s��_&[�?���Z��I�&4�h��Y�I�h~�:��d3�^�Q����"9q�Gș�!�j�a�x9�e"��'��Q� �C����
��p|-5��c�qWMz���+�n qs�m	�9e��:��Ӧ�A⍊��U�h�2�(��G�[I&h�<-[��]�j�<��Y�AC_�_D7�s
p��yd6*^�]b�|�O�>�����	��!T|����sN�p��z����^�J�x>�Gg��J&���:�6�Q�t\�A���p�U��	j�������%K��&�}�gf����ײA���s���Dq/ۛ<�U14����CĀ=9x��Ѵ�g�!q�RO&�v5�i`�"��2�N*fx�O�W��f�[�JL���t�)}9�a��8Nժ8I�ă�}�>����� �5�R#�ٔ���rg)�����@l���U������=��)Pt;�6�	`�1=����9�-~��X�kP#,�}�l"P�vk8�rl!h��ܶm����|q��
B4I�˵�T����7���-n�z��VG�}�ڜl�,���v�z<�����?p�t��b*b���$��׊�L�R'P=�,)S�"�L�"�G�WG+��:�� �Cm�0�}D���2{^
4Q'�c����U���;�//���B�ZU%7G�N���yu�ݥ�~7�7��R_��7��^��Z�G��8D�ʙk��.e�� ���p;=���l��9����QŮř)�x (��~�HG|Ω>��Q�e��NЛ�s]�|� rl���&B���D��P�!���.x���l'8�OG���O�V��s#�����uQ������c�@�M�������p:�-�|����b�܃[���KM�AW�t���v=�\��J��K=�هPS;�h�x����fsQ�����r��k����p/l�/�eE�o�ŀ��zn!s]+?:+C�p�����ǒ���h7e�	5��_C�ʌ''�'a0e>co&�Y!"ǟ��ܠK[:�.pR�A��F�*hv��
��'{�%j��.��� a�u�N��kW�C_[5�L|�.�1(	W���DL�۝�c�˶�a�`�)wuhTmv!b��@)ao��<�ܯ����r�[e�Mg���6W~��4}���,��Bq�V��1�kup��\S�ٹ(�����d*�^D�O�s��C�ord1�/��(}&��2�^^���Tm(B7�Q�!�8���6�mIm}�YuF�2����t�x7���f�Y�q������~��RR�+��-	�����[����'D�E��2���_?�[aKN^��_PK   ۍ�X~��k�6 4 /   images/663b53f5-e86a-4272-a51e-f5b809259b46.png�yTS��6D��U0�*�n�4JTP��� ݠТ�
A	CP�y��j��mQ�L�4�@ ����@E� 4$"B� ���пw}�ߟ�ֻ����^<U�k�g?��u��/������[��O$'nE%���W��o��� ~,=󟟏|F�W>𿿦�t����G�ɩ#��/ׇڸ����;�7:D;s���(��_��b�	�3��G"2G))�)	�-�H��[_Ɨ�e|_Ɨ�e|_Ɨ�e|_Ɨ��H�<�/p�������/���2��/���2��/���2��/����bl�9�Ϸ �?��7��S�9gζ���Mт��řv�����'�6~�t�y뽇N�ugKZ����������E?�G�'���O�0^}b�r/��̪�=9�����g4K�?E�d06:�b՚*������2��/���2��/����6�!7������CSoo�Q�ا>�:��3�"�ܾ�yT�_Ƴ��1\�yk8�v~�V�����g���d)N�.�х�I�3L&�}z��U�B����I����Os���:�O�@�bt����j�A��,��YZ�Qr�p��`���5��^Jt�l��3g��g0�������ҀŌ��~~�hcG����a{	|�K� ZZ��,��%�o17�����2`�`�~r�p�*3�������(�w�2"Ɂ���@�hy��ON�����x�*���/lU��b���].�?W�-�H$+
?����%{�1��x�EF��*�2��K����AZ�� ߸�����4@��_0+��r�� ���g��O���D����N�ʲ��\�C����6t2*�vnȺ_`�",������Y�;����Ui-j����L72{=��H�5����CB�:�F;���k*�3{vaa�q5���[X@���n�2T7Nah���-$NTײ�ڐ�����	]�8�scO�*�XwF��)(7�x��xλ��r�	�F��(��s�����1�QP�Ƞ~���4*��M<7p�'��Q�A�����"�t�A���t���#ڇ����l4}����c�v����b�|bTx��DǑ=���M&BI�$������.�k��>Ը|�B���C��VQ	Z���L:gO�]9����C'�K�Q�x��ߵ?^˫�S��ai6Ǘj��:ٗ�`4|x��Ǐ�_�~��*Z�&c'ո����L.����\쓷RE���a���<�g�$ݽ��̈�r�3'�0J�����:=�3#��a+�^�V��65�Lm4�����Ne��w�7S3�9�70^0�͈����Y��K(��34=A�)WB�ێ����%`	c�y��j^�1��!���Rc�	1�'��p�<�M[`L ~��*3���gϞ�~zi�����'��&�\f�1#��4�j����]IG���C�������<^ֹn̎�1;�CvOm4��bD������:����xY9_"�ğ{t{[!��9�	�9�^��I�s7��'�b<IT��V��1 �y��lb�H
�O��ƞٍ�݄(�S@���<H����$��Q���������*�� jA2�Zf9X_c��i/Gӵ�����={6(���������	�#���Tr{��@y�?~�O>����~c/o����J\��ê�Ȼ��sQ�T�&��`j�11�<�C��,��
NW�M��}�*��<�~UhNHLө�����N/M|z�u�~zԳ@��}�<9����>b�F4����eЈ��Ӎ��֧6��0��D�z���j�4 'O��
TL&^rd��z�s��?�iV�c���4˼��i�����^�� w,>�qt=��c�H�����¦�F�������To�z�b�!~ԅN�m��m���NAn�>13��wSEB���H�zE�^`M��F����W +6fo��I(ƽñ�5�!L�~q�"�qP�ܞ̜��g�A��m��+*��-��f����-t�3�B�u�9��`����5����h������;�s�F�,���Ը���3��G_LY�f6 |G�����#��n#�[K�Dp6�x��}�o�=�{��x=��b��r8�r'6�̉������.�\��]��wz�;Ñ��fG��l������mG��C6�$�'��]���drd��ߘ�F�/�M&&�3�/|N�^���7xօP=\�ۭ�
2�hƩ�VS%�w��>t7�ޓ�lu�;���+Qm�YP�����D7y�s^N+/����{G_�\��F����x�|vv6���	e������?lf�J�����ߧ3���_��- �:�~>�fE�Bp�:�|G7ӬEIĕ�@s�&9��ͼ
Q33҃t�b�\v��=��7f��Q�n�C~��^��ӯ`K����4d|c�3�p���2�����|+3���MhN�+v�՝==D恾_��.6��3p	��w�t��(�EE �B V`��Z������-_8��w4ՓL�VJ��gLSɱ�eq�.E/�v.Ϊӛ`j��������]���	A�u�ݾW�jS}RwCu]7/���E##v##��-���x�'w��}M�������r�E|+��Ң�����A�@Ɋ\�Ew�{��]G�p���̙d�a�t��,m�_Ѵ�����������_w�F/�PW0���Idjw/�/��0_:���}��9)�s�
?t���qt:�SS`U�jh�����]��?�ÀBj:�'��/0�����q�<쌮7'Zs��u/�jF�>�U�,�T�;�O��E�t"�qF���o0s(G�FzQ���jpئ�sY�c��'�A��)fNkK*�}���ݶ���ej�W���p:0�
n�I��,��،`T�QR��W^^�>5�9���=��*��U�쩔��mD� �y��z�E)�lA��i��v07��r�m+������X4�;� ��?�ɖZ��הhiSS��%�%X�C,���:\QΏ�$,���.������?�.*�*~XW'�KVw�1���s��C�J���|ud3���F9��{��̈�EZ��B9�If����O���0�O��K�B�W��6Y/�>��X�[���]X�|a�{����x{ژ��~-��b����@W-��z6��
a׾b7A��=m ��g�26����6�K	�bq�H�	D�	��6�dE��=���f��0��܍�!뺺�ɽ�F�������_��Ved�%��<��陙>��"
0v�:b�(Z� �F�����cG 2T�ysA��0-�Z֙�O�U�Db��L]��,�Ί�֫�����J���+B��&��>�e�Y�X����<��s��y�,����r3T����H��ŵ-�ڋ����y���ڨ�eO�Cql��G�a�/cz�f�l������~�����ݻwS�b��,d��n���0Am�:�R 1���L�".?Ƣ����w�j��橐�]������+d��b/�S��E�JlA&R=F]8M*�.�Y?=�}~W��ѣ3��l�t��[ I:_��,���S�NBG��S���Y���"��o�E/ߙ�eJ&��#�1�% �0�t%C��y�n� �G�Z�="��K���LФ����?���;�`:H���pc(J��)�`��bL��ئ�ZW�c(G��`%驲v��j.ڵ��������B��@>���k���\�7�,�h��յA��{\56P�O@Z�'��!�Ȭ�@r{��H
ڷ�K)�!�L�� �;d�f�i#u�M��y?���A-���,���W!��x ��Y��ߤ"Ux[�'(̌�y��Wi�L�DD�u"##�o�R����N���"��&�����?�ݎF�"��p�U�6�E���"%���u�s{}�C��oѳ�A�����踙�7�C8�VO&B=Ȗk�Ҭ��o2�3Jk)�m�k!(�̒Tn��h=K��L�6a�X��Dn��)参��9}���Hr�2�b#"h#���
���Y�bՁ�G�g�uT"���+��Z��U� ?7rX4y������<�vP����u��$�F�ҙ�.�71��
JH����}9 #6�'�@'�tHc�B��Ħ�>:@��xB@��fjY�?A؁��M�ΉN�aY"6W����1N�����=t�����{�Cn4d'Q^���Rۋ�b����Ug�ꔵ����������[�V~���s�1���Z���⩑�S~���'ZZ��+�TFo��O;�pZK�J�$q��Q����U�j�0Ys�I���D�\*sfpp|Z�p�Q��%5Һ�3n���?�Ŝ��{�����n�1;�T���0,Tl�Į���.��oMd��%Q`���ۉ
��빯Gd�FL���=�O��+D������C�y�`��>���D���M65�&ƠV�3��_&g�2����E����A~q�_��j}ʹ�vR(�ܿFP~f�U7w��G��%ݩ�w���J�2]�z��`���-TN�-^=�葆�R��Ϯ�K�7:5Ǧ�58v2/f������\w[f���vl ժ�?+ ��M��U_a��@�y��TF]P�J}��</�o�d�(b�'��Ю�yi��k����t�RI���<x@�bo�w4R�i�z@���t/L,�l��Ż�E��9��#�P$̔�r�����n��D;}6z�:�aC]��r����^�� �ÿ3��:GA���������0p4�A����/>�=OKcv��'Y��>=G��:'XO�}܅y���k02^�-�>�T:�z����~4RN��蚾=�=�x���\��s�����4����ⲟ�u�\kc��e�X��&L�a�_ �[�sl<M�u�yٓ�,�S\��Y�41ܪpk�	ޖ(j�������"ń��>��xG(S<��]$��s���T�؄���o��?���~sÃ�#��= ��E�@�����Қ��b��Ӝtz!b����t!�N����ǟE�ȟNv��������� ��.���ZW]z" 5Z�~i��co��5�b���ͫ�q�y�[	����R���%F�b.�|	9��k/�&.����������Q
�ѧ?1��g}䝍�&̘(R�-i�s����5��W���'���X<��1x��_��'DNM@��tu�u��#�W��a	��������P�34އ�`�'��R��I��!�ꆔ��쓁��t�jl$���"6_k��xqRV`6���l�p��Ю+ Qe� tW˿yr���!�/���'5��c�ׂ�4J� �S��G��#��7�D͑�>���`]o=�,�t�9��=R&�MC/ӭ÷k�rѓglb�jV�Ps7��t��1��rF����A�%\��9:�}����g.>ygo��E���|����n��ٟ�~�QP�4,`	y��7)b�[Jpq���1>��V��,+��w�^�l[�e��,�U!�4�p��l�쪍y�-^y{�9oP�E�f�o���*����͆���|���^���X$�^�e������`M�K�x|,���s�}�Y�T�Z|�~��_.�)�j�̴bī1�E�
zvG������`�\�t���Fz��s6��0b��5��9���~�_o���	���?�h�K��T���k����կ��śĀ`BZ���Ț"��wQl[x���	gM~�T��&�͗�6��[+�	}��&�Հa����0�K��=PP*��0^z�n?����S(���1So5S�Y��E���˜I	��avS蒶��ܓ�/<D�����#�eޙ��
M6$�m'�c��݋9�gw�e^ڧ�:5ma��o������b~v�C�{�W}}����JK�UY�
�Jc�yccc����<U���E���9YL��Ւ���wA�e����Ë=�E�����*	��XY2P) ��-��t)8aKj����ж�*�vk�dS��XZ�@�x�SSr����D��Z���,�x�M�}*;�0p��iqjʥ��o�y1� ��G$#��N�d�zK�2�}(��?�|�u�V9�'A��1B�nG6���kD��c[ݎ��Ps#i�b� W ��->M�,?�'�!�� j�a�[�`�8� B�8��W�/j6��%�C���b���mܟ�:�B{�����������MaA��Cq	�k�
���&h(%p��a��AXR��~dM&�h��uR�������,sٻE�H:
��GDߛ*g:�	�_��[7�&1l��u]�W�2&�MXo�u [ �p����d�Y�C�d>��w2����@+(��T�2�#�@ �)cF�#,0 �^�K���5�j�D"����;U��� Egȏh��}��B�t%}����G��27"�0�(���I%�:�8wGd�fUUպ?���6�8�Js�
��)���-�@�ʟ�G�ز&�~T�C3��^��suc�4�]�ɖ�Ѥ{�"@|3��Q�&�~^o�l����x��%D#Gag��n'�@P
#���u
����b� ?���(���13�~K������6LH^�o���"�Vh��c��?����#5�QNiڧ�NM��JwJ��Z�#�񿃏�7��𨋙����.� �l�=�")ox­�$s�����4�Q�t�0����c(��dJuT/�tCI�Z�kP����my���E7����zz�kC��߀~3��>t�ҩI�� ĸ����T{�z$~�*�z���4ˡ��?�٩�,�w���h�m��B
�����g��]Cc�YT#,�f�L����"�<\b�h�͟�+�5MihWTG�am���E�i���a�B�O:	�˹��y?�dc�a�"�Ƙ�,�����&���d
�Ks�i�@��v!��6�Pq!9T��3�U�U�Y��j���L��2�o�1�ڊ�[z@��������S������lz怒���y�!����������#�v��)�A7��ߓl��[�;=��Dy�d�`����@�W�|�!��a%�H��+ȉ�m�'t��1��0�	4��E�^���l���#̾�ݖ#���yaA+]�ۿ���O����a˶�㫀�ܹ�Ҕ�P���7�U��U�����P6�#w��'J�kC7�a|�Z��XS��A�	:�'�9�*'^<31,��;�NV��2#� t��;O���QpA��%q�'2��<g@�b��G/˴uu�� �]Z<�������
�=|��`]W���l]|{�E�	�V�d+��Uw�r��x6�-��h�����*uтj�j\O4�ßMrjrFHJXr�xX�F<�A`K�P�x����ȯ����T,_��Xm�N
Z�Dr�o릱����cݘk�%��E ��:�fek���N\$ ��ҋ{+2^(kݘڨ����	j&�\_t�vJ�Q�@ģ�v�z	Q�$�
�}�Oj*C@�pC�`Ț�'�{��k:<��q��&�$����;�����޽�c��S�T.dB�2�`�����o(ZR5�Ӈ��ݮ:�H$���X�y����j�T��wj
����.徙}���kTAY��TU8����WKKK�� ֗�|9.��t�ZR�e���D j䥁�2ѩ���8�{��p��I��kv� g{�`�l�%H� ���NfjѠq�:�s��]�{m����p�3�����N;��*�%�����1��;[4zT\fJ&��re<����^܍�CB�5t?����.]r���BI8H�i�4�P�W�(�|�3�`���N]��� !�v����q��<
�?����QX��k�G)�M����ԖO���c�K�k������I.FU��=�YG_��kD���k��n�����
�ljh��&dHۛ�#
��֎m�rA�Am�`~�a`&/�$����bs�����0��˥��6��l�!�1V�� Oͱ̥��#e�����\w��A�1��҈�ҋ�|�����K���_'�E��sCﷀBQ}�\�����I�?k�&/�v��Bv�M��2[R���~mo����z���sf˨L+4ӎ�
�k1�J�hٺ�=]�!�
�Y�����N�ꦢ���0���6�BG�)ׄ6��Kq�& :s��U�#zĝ�țnD��k���{$���}���y:�>,&fn���$b�3�F�T�f6?�������N8^ָ�$B�5(�d��c��g�C�����߂�V��
3'���g�U���O^gm5���@��x��#����_��Pƿ�u`���_	���������Qua�G�0��x�������	� ��)0������{ī�o)9��n]@ݮ�������ӸX21Pm��
H8V:���a��|�ۀSl�)�a��`�
3%�S���'^+�4nq��
W�T%@�m�;7�$#͗`��N`fa1w�C��3�/���%�����P)�झ���	[�]^ܾ���ۋF����ə���t������@����)߿Mw�(g�f{���z��1�~|�H��?�鬈���@���V�܎p�}�?4�3je���^�^��y��pKl%���HΝD��ô�(������myl��2�Uf�sޠSS�Tn#ޜ���>��w%��T���aq�0�P�kk���s�څ[	�91?k�]��Y^��nV��s���Vtm���js{����8�yF����ů�˃������X�����X��E�#f4�Yp���r���\�|��&��/ �S��Ry�~`�R�q���tJVVV&��O��0Ǭ״HGGk����0%�#��VRr�=����$8�mĉ,aW����)�y������W./�/ȁo�`Q�f��,��`&32�	go"�?p�y��V�L`ַ� _8L�rCP��C����U���V�N0����C��D����w��(o�.�l�"rL{[���B��NI�J���"�q�S]�s��G��=�(�yi��7a���B�N�6d�ks�����a����;��C��oa�\<���O��s�7n9!��qV�����P]X:R�)v�����
jY��?˱�@�Mxq]��mp�J� ��L���f�2p7�1\�ূY����tY�OX�@/{
uKEJ��^itgo�v��X����3� ��""t�N9���.���A�~O�p:ل8���(�e| ��h<9�"8��B��M`������CuP~�_���/�����N�֟�V~�}(�KuS����)M�Ť���Ϡo��@�Qx��7�"Vux
j�Cq��uW��x^'�k��l��u���k�l�?��������S L[z�@��;!�]J��)��"E'w�����0x�]��kCE��r�vAX盛�o�?��O P��5���D�p��	a�O�0�9B�� �T��iM�|���[��Wl��5�ƌӉo�D�@���)�խ�	Mt����9�u�E���yi��Ņ��V'>=0���#��!�T�5sZr���������mE���C\���w^�K��x'l%w�t�SS�u�Xf`�~��1E\f���si6�N�G�>jTNT�6��ۧ�po��jGGGb����Adsj"�$z:��{�B��r��>���a<�e�$����p���x��s5����!�9���0m�5�.2�%�z�� Z���Pu��})J��̙x����˰:���W��᥽~ry�_�aY��zJ�"�;dj�i�g��Lk����Tï��A��&۟V�k��=��mi�	�N���;�w�Z��J�sv��ّj�>~�����Y#���{���|j�>�������a�UNv�������q���+�ԸO^���>{�uC�#	�@����N�n���<L��V������e�,����ss�P(�va��֜��'�H�/ Y,����E�/��+�^�v�C�<�mꉹ@2���+]�"��~�KP�5hs�,�/ZlUev�=�����i+�^%�G��}���pa/���Ga�	H��d7S���^�0���d�졉U�v^Vq�`m叫A骏�Щ����(��9g��ʾLf*���R��TH��I$�(��2[��G��:E;�+E��X�O����ɰg,,�����#D��{K��;��B��,�Y4� ����ҴO���R�Tr��a`A��Z	�Kg'\z�^�4�;�,ςb�n��VB5�Q��f�'�0��������^�ϊ��	½��˲r��i*�Z*�s�;
�������U�X��:N�����J.�	�Jm�ވ��E���cK�78�Uw���s*T�*/4B� �_����?`%�׮,���P��o�\���}���G�`~��2} V.�;֠7��~t/��p��f�"�����;v�\~�ͯ���#ĉ�\��;�\~㑮,V�p<b�6ݏU�
v�:��\̮��Y��u�#���Lv�	t�?�</�8lM��aZ,�9��1j,�l�MƁ��cՒS��U`9�H6���|(IP���;*�5��%$��䍃���.���Jl���0`���E����e���!$&8�z^���	O!Z��C:t�=z�(����Ϙ�8�"�`p�����ea+K#�������כ���T&�T�[���L&�771uRyn����+���	����l�p�n�j@#:7�w.�ڝ�K��-����S��4!J�aKH��������?f�1����cR�J�tz�,|�+��lq �l(�W��[�W*NwLaThkiYTayv��d�e_l|���,�ͯ^��ޢ�@�ZW�H7r'K��t7&�/��.}�؍#T��@P�,�С'�Ń6������R�g�d�����u�}������5���.���m�Ɲ�qb^Z
�{0���B��}E!��]�����'��)#�ʷ�^��a�6d��ϗtvuE����<�q�����U�1#��
[���R�u�]��
A:����sNPpp�]Ҍ�0�w�lMq7h%�)J|������w�ޥco*7@7��ߛbq�f�kXCԱ^J��֨Z�o3!�d�)P},,�ſ����x�yԯ�3ն�]˹����]Hk>1��y���9V�8h������a��L�̨�Y����8l�	��Y��oD�K*��P���}���)֟ڮ9�ȘNB���(�N�^i�����7CL����J��$��맢^�4ɟ�Aʤ�*�?���@o�E��/�͊˞<yR��+�ӿ��~G\���������_cƿ�����j��CR��_�`'�k��G�w�<�W*�Y�
���﫽�]��@��?�n��n�0�4�C����Za�e̪��8{�W`� ���/���(ͩ/n��P�b�[�}��k�|-��C��e�c��6H�!�,��Ĳ�^墢H��X(M�%�����MΈGFFV奕�;���=���X�IX��a���6d���;��w#��1[�V��<k+��M�',��{	�v����?�p��U )�@Juφ�:6�
z���huê��| �*(0pޝ�[��{/�ĿW�p3a�N����0�fjj��p�5J���vg�z����k US�Τ�rI�:���ψ*���D���j���+�1�d@\��=��Z�=v]�b+�}�?�k�H+3[_��`(t��ѹC(�ϼ�X������ٻ�{��L�r>�ty5�c�:��������Pيtc��TT�"(
̖�|�;5�֍��"ƹ�艫�*�ހ�u~|�}zL���7q�g\mgF��ޱ�@�3,R'j��Y`� ��,Gk�-o:oi��m�re������-?�����o�D6�]��tn��/����t��i�b�#,��`��B~�X����4�)J���[�e]��|�f[�4������F�@~�B�ʍB�cV���~�Nw�+B�zwd�!R��0����_�f����/������k#Bd�6�i��#��v��x[Ľ��}����M&��ߢ/&\�!0\�u��
o0s�Ql�� SѴ�26CJ��J-�(�p��wnH�^��[	gg~)ĀN���Q��?o��b�|�v�e��n0����k|E�����o8��י��h�; W-?�kY�]�3���v��|�����N���p/A�%O�0���^�Yi���5T�_�4�W� sY![U�xO����9Ō/�>Ü9@��7Њ9���2`��v� �����E��y�o�7H����?�d���[��`�G��������: ��1xZ�;)I������b8W5�dW����L�#���TE������<iψIg��w�Z�R� ��>?2���!O�o���3��d����+�
�T��� �YX� �k5��Y����eh�%8��e�L��^�8U�[����RΗ඗;�F�,�DK=�K�����SӇu{�(�W=;���;7p�f(��ynk�_��<�����9�+���flHI5��.4�)J�6�4da����u�rww�K��,//�
���]q��U�dQ���Nv�q4c뀱�Э��"��7���w7�S���C��A�f������8���#9̒@�`�mh 魗��-t���E�=�ܜb�7����)���=�'�'��&�_~%t(�����l|4�5�;mm����K��p�E��_eÝs0�:�Ւ��Y�r�䮝�j��������Ty��͗��K�ށ���Sg\i�O��G�s"�E��Xa��Z�e8�u3�n��@G�^�I N����*>��蚷�1Q�FLݝ��%CVs���'&e6����oT���cSb勳� Mg��6y8/�Uf�,���J,K��ݨ�jY�z�%E�Ӟ��;�%A7dv3MfUG�ni*#�
CԚϏڀ�x���b�����	���p��]����m��_�pt�&�j�L'c:9RND�I�L`l;��Ҷ�e���Z%9S8/�?��j��}�Z�H@Yg�*�G�<��?ȗ���b7����-�O.3��JB"b�U�~Sj�����<s�ڸҍ�6]�Rŵ�ɾ{�l�>w_¥��x����P}a�4��WZ�3��TB5$AF��W>�3��l�ݱwi�&~<Z ���EW.'�o;����4��g��d��j�p�����HV"[fff���/�aG�-��ɩ�ʉ�#�Sf�5���O��r-�{���t:T�.]X��R�b���?��΋�nooW���5�̜ P�τ�lT=������~E���*��1�`�ҟP�^7������g�����\�!-�{�o�ӷ�5O��8JZ��e>Zo�Ӫ�ԃ6����te9��B��tj*�B`zr��c�0>��}�ǻ��sL:?8�����u/������d	Ď�z�X�;�������^g>����춾Ɯx�����\5\�)c��7� ��������G�U`�
-��zVR�Oh+).��M�@.L�#�MLLT���*���"@o?@�ܻ�����V�����ϧ2�E��H�I��;��G}D����C�Њ����o�g�y�&�*I�*,rZ�	sI�ύt`�>��Ϟm��[o8YE! �SR	�*�׃��/y� v�2�`[�ƚ��$��(p�7?\�ɾ`���3-֝6y]��Zځ\c�8/������F�zJ��c0�N�,�{�z��2�Q�0�q���Tؓ�G:����Oܜ��k�8�@K����h/��bL�ē�[�me�0��}RJ`���-���sQѹ�Oݺ{*T�t^t5�T|zJRj��ʉ,sb?��T׽_綍(ܛ�j���L�kH���T*;�6S�l���#��[b$ ��I)0��ውR�?9(Kw�
B��T>�L���?�S v���k��I�TlbjF8P�4��v��14�����[v���+��k���8��R����P��_���h4�#i�9���IW�&�N�Ɗ"▛�"�<��HO.M�k�ԉG��I���=,�TD���n�Y�G&~��;񂗳��j�-~s��?���7�'���7��8�Y7P��h�,�K6�%�%��D�C��O`��L!��6��d���V��8����B��8��򪢰�b�i�i�L&N�u�$�a62#�`��N�i���7�G���]� ���؇\&0����_�ϱ�^������������}5kzΙ_g��� ���Wق�}U��f�.܋�p"�w��y��P�~ۦ�g}_g��n�����&�m���~��>L DK3�� m>0!��Gw�%�_sV3��u�P�l�ٟ��ͷ�x�,v�GV:�{"'櫞�T7Z���D���^T�'�Ɨ�V>�,�/��2AD���¬2�{�rPf��e���bn�j���F9Gic!�ɓ��o�ic��,g/KD��E��@�q��� �8ƾ�g�\-�Me��TV(���v�Ut�Cj�c�Q�H��O���'�V�*3#���+��W�:��Y������jX:�[��p}��e����\+L��vL�ǡ���-[c����@A��2؍0@$R{�">AҲ�Z��r�e���"��/b@���`���q3��骹@�e��w��2�����l���.�y2��S������A�,�m��ڗ�S���'e��Axl��C{��kim���~�ʪ帞���3C,v��S ���0��!I����:�����P� ���%1�n�͕D<�-�SZ�"߫f�����GQ[l+p�)|��~O�.���O:��i?�H��fP+���O~���2น�����+��[[#��2��F���'vgpJ�N��"���<|D��Y��(��5W|�6AC���!tSu�5|�+'<�����6H���tϨ������Y��?��:8�d���={e���� ����]H�W曈�! c�J~�mՌ�ԕ]l>�߸�#�	.��]!$��wǂ�"������@�iY��j��c]e�!�<<�u8~��~x�"Z
d�C�,�l��J�6T w��WrҜ �U.W�E�����:�x%E-���z��{��S��G�3�hN|:�g��Tk�:�)�♿w���Z��f	�$�S�N�qhW�v�Ŧ�͡��o��mx�.!Q���������8�
������{���w�Oj��'���T�9�B�����E�:��/�{g�i}�g�/��?m|�	�əŶ�����Gc5��˟7��k��=s��6�.���w�lK���V���C�(H���K~i2�������V�ϯ��zy�'o�jw���<�P�TP"[���u �;8�Z;�::T�G�[~Wyv����9�ف_�p	т�;����W�H��p%�G����Q���EPAZ��o�j�*�B�x��Iw*�z;%X���a���M�b^j ���S�E8��L�d��%ĊD�����sX���k𻀄��1<d�'��=3�A�#�z����j>k��{$)Fh+X3�_Ce��]��AM@z���<B�xKI�Xx�#"Kc��pޠ="���CWr7^f�r�&�\ ��;�z�IX�D�ajn�t��(��E��#z=�����w��Q���KX
���o)n���4˦����ꭻ��y��JV<E4ō���9l�-����TVN����>j�hH���{���A���Q�Ұ�Z�!��Ȑbj\v�ۚD�r�=���.3ŕ>~��Ȇ����+�}���bhc��(�7��Nu����F��yP����%��,��ІDE������D���L���P�U`�6Mc�UW�oZ��̢B/��i3�qX./Mx�Υ�ƶḌ���ڦɝ_T����i���g���$\�_��h|aڧ)�?�g��95��M�8�T����>B�Cj a�;~�)���}�Z��d���Q#�i�FmX�jZ�#@�����츖��R_Pz/�P�T@~�H�Ix�a�?��X$�Kj�Mg���ڵk�:15<a a9a t���w�QՉ�Sjg̏Tn =��֞vmM#�_�����_��`/aLL�\8���Ӄ`��@���9�Ņ����Ye�mO�l*�]x�'oQ��<��-4�ľ��ե���)7@#��/v��⒒z���h<����������k^Y��bM�5=VcE�&�֒o��"��N�`��?���H������m��2C|�n���Ë�\���̳iP��~-/�w9纕��<�f�.��OdP e�=�7���~��KSD[���1×�\c�r��f�;5�Q�V E���w�b�j%/�Q��/?}�O6p��_Ɇ4�gʑM����ƛ��,�ih�^�u���/�T�qP�=�fց�丸����:G~�Ƥ)/�%��e�4TϏKu^!�ѼKW-���<���2m��ψwL�)�������,�����=�V�$�E��΃�m;��Dw53���ܝa�CA��������wj����ȇ���	]QZO �������3#_�N��w��7�a�z]����	�ࠠ��ϟ?����	��)��j���$��U-��AmJ|���m�G��,�p�#kr�����ˁ%ʝ���lA�+$;ʡJ�*�����ǟQ1O�Y��L�؍�5�9^>"�H����0�\t讃miǿ}V��g	!l%-���5-��[@v�������*���g)���,1�(��i�d =�(�{v���DJ,��A��׹���Px�gڨԏ���{�[����h�]�俈��~c�ɩ����="ԟrb�%���QH�����V�z ��c&g���FFF}!@Ӵ�],�w�"�]R�y�L�a�;�p�'�Hq�����Ι��k�����&挱z�S��� n3 0�G�	�0Y��6�DćPb�O˼��N��ߖ��u��	"|����s��O?�	r���<=>~	S
�C� �� �XA��"q�B-�HR��΀��چ���
���}%wOE�ӟ�L�j?�1��[4;��2P�kl�ŀ�HP��G�̙`�DSvPÂ�h�Tא�=�I	Xnj��{y|D�'yflW�8Zs��R�.HA�|�yN+(e6��h*���(��d]c��]j������� �'���S}e5CB��S�� g��eM�w��A�i	cM�_���3wB�5����:D����Y뫕[�KJl/qo_f�[lK��̜�An�|�in�(�Q~�c��f9m������O�+�G�Z	o"c��"�[�tPkY�L�U}f�4	,���:˒�Yb�OXp�<$k���2�;}Q�>@�PjR���}[��~^r��Y~�΃�Nv)��'���~��{���u�3���8�0�h�2�oÚ<2_zؤ�Oi�����SuV޺;��5�;����3��e�+�>�5��3�.:Z�t��%���Dqgg���Ҏ��j9���,~�^ ZDI%�37�|�_��|L ]s��Q}$�}I��U�O�7)�݈��p3�����A�wD$T����`���T*綽gFvF��|�DFKK�Bb툟 �KmA���`�,>+̓�/ׁc-���C��^��w����?M�^���0�Ը!��[P��[����ڹ;�S�yi�I�8��;��� [��CPF�u[��������aP.-S}���4fnz�5��K��]��s�������f���ڐX��u�/Fk�@qBz
�]�`lV�n�m�:�[f(��ù�����\���]0��~^�37"
�@���ן�΀U2�⮫u%@�^ P���'1hEl��o�%�$�6T��YBQ{*�Ea�Y�������{ a���npj�	��넷�/5��)�[�z�$J�}�lQ��L!�}���ߨu��J63ǢZ��g6{�^�i���~'��N�:�]����'���o�U`�{���l�����qcO�>�݀.�e/N}�+�¹B@���6�?J�T7��y�* ��\hY
�Ö~�E�#��1L,������2*� 2�d������@�07Hf-KҜ��Bم��f�T��^�� ��|���i�����l\dkɭ��p�'�Z%@�m"��|�`�?������h@\PAr�@kX'�򧥋��*LrZ��If���8���J��L.���I�S��Y7����#:?�:�ɬ[�4�&/	^9j��S�8�L�`�A<���eI�� T��C��ޔ�����<�}]ϼ�ނ��m+ùw�7��S�X���a�(���b�[a�N���h������i��H��"�� �ςh��
�a��������5�@,Ő��ݥ����Rw#ŏ�1cu�|%��ږ��'|��H>���л`�X������MP��5~ĝ�q���[A�*��	8�6xA:5���������u�����o�:{�K�ڊ�m7�\j�]��!�]%���P2��Kr�M��"�M�vkQ4(M���&]�&+CaL��eH	�眷�����k��s��<���������Ґ��K��M�$��Aw���i{b����`��@-���q$�kq�e!�b���6��4���t�������_�ΗFVg"6S�װ~Ov�hY��?�a/@�|���LFM!$³�#��˿#����332���o� $ j�L�{�!�z��"S3H�T�K_.L�
�vg��;V�Ul�{�\Cgv��!�z$��Xŷ���⮐�v�+V�&�v���u��V�V�N�{r~� �x
hPKR4cC���Ɉz
������Q'�G��J_+4A�\V�e�ҹ��D;w������OY����@jF�~aKw���
�X�R?/T�XH3�5���L$�#�(R�=�.q�?
P�_�&�2�a]Q��(RH�03�~V�{��6����� 矠����I��|�X��Xо��d&/��lc���ެ'LG�%��z�y�����W[�S�rj�{F|�o�W7|��jii�-�;��G�9�@Y^R��yx���Cg�f�#��:O3��kb��H�m�`Ψ����u�1��9���(��npKV�+c`��I�*�\.ٓ'���[����S��D���H��#`:=6?ڕ��d���.6����H�$�4<�m���7�t�,��W-7�����TA�7��i%e���[�6Az�J�V�t|F�	-:��R0�$�(�&S�*�B5p�5��[x� %��|�C�K���z%s�
��0{RZW���Y���k�S��@�y�͠��!�'�%�b���}�m׸���߂k��sZ	�
�~�ȓR���G�TQ�x�/n��,YJ����;�DZ�h}}����:�t�U��ji��_��%xÆ�����hZ�B�mj�]�h�U��r�^䠘��2z��|����Ѫ�����j�d_�n����WK�}�����'a*��E	��9���VVU���}�#(nK��"5�`Ah�U��o���1/�������"�I��}�T��8A�%�ۨ���|e���%��oq6��|l%��+ӆ��ž|�޺�њ'L�F��7���S��[X)GӤ��ܲ;��:���m�L�t?b"l����7MWԉu�0��}���gtRx��ѵ=+Ge���po
Z�D }w5���q����� [:����?��#t�755��:U��->���t���1���dYXm�D����|�� ֢��nk4�@�8��Ldk���N���V��N�����:��H��=NdU
{�A� �Lu�|ŋ��������>�>��Q��.1����;�z�Dښځ��+����+#��y�5��<0߰�H�ڹ�xT���ka�ͧ=�rU-C�1��.���]Ƙ����#��sd� ����<JC)���v��5��c,�f������S�tDai���?dS+��-�'����ԉ�R��r�e�"4*�����G7�� st�o�#4�揦��U�]�wS���(�ܻ� VTGQ�ea��OeБ��?���`�Q��8Zc3�{\��1p�_�U�)�	Y�*���:F��}��)���IB��Y�����ƶ�����@*�Q��W���Z�T�_�xa:���g�)���mu+�%��@�;A�c�͆�;xo���b���c|��96
�(m
la��2ާ���)�@�S�������Ĝ�5-�ãr;�ܟ?8��2����^a@�ru~s��0;���ի��H��L�	�'@����&�FcZ*�詶	].���,Sr�:k�>���s�S�`z';�Wbb":�YA� 2�����ʗ(qgqF�́E�h�N69�ri��P93���[�/��BW�@L:�Zj_�^E��o�X�ʅ���V#�Ɠ�y�+E�A�Z��c��^o�=߰��XA`vbD=��%0�:%�S_���gl�]� \W�ŕ��J]�ڶlҦv���u��C���ZrBT��=w�0����۫]�\H����#,���GO.(1�����C�	iM1�jM���9��9�w_\���a0��Ӗ��Hti�.v4�b������#b�I����>wa�貈��w����[Fi��OO:�wQ(-�����.�*�p[�fϘ�?B�4-�]�-#��a��s^��dGVEch�>�
(���W@�q�L���]!a;x�P捊3Q���x��&sK-�Xl>g>5���p[�ߪ�Ӡ���ʋN���TQַ�0�3\�o^6�Y��YI�#DQQ�#A�ԁ�(3�zmkFq1`,i	 ���%9�F~q[��Őa�����Y �� �y��ǧ�b@Υ�;ܣ������Z�����7�0H��iK�OP�Z�	2Qr�in��~(�w��k���K�09re��f���.9�$d���H��ɱ�'Ն~w�y�V��.H'�Y	�G!�wzݗ?��5���������T��/%W�S��TPi6��'�T'���F��݅���#�	�_Q�ָ�xi��Ps�W��h@�)�{h�whm���zuJ���ܬ�0�]^c��9�o��]?��i�~� %3 ����v�2��I>Ƹgl鷪��g��(VL�Ku�_��Ϯ�M��T�zFa�
Q��hP ����ɗ��g3���mlfڰ��W3�!����c�gT��H���Ooo�x��AȾc���b-��7.H+O.v,���N��㪻h0�ka�Ç�>�����y�FUP���u���В;�!�N�.�
�T:���	����8�u@E��db�¸XWGgj@��N�U����;)e:�u�8��oe�wW,;u���Ө1���
�)��0���7���%�";J��,�,�6���
�x�A&C1�n�I/�0?�mGt�:d�a���V酉���]�[M��Y���y�>�)c����s?��F�+��V49��a���w$V�j�Z���5\�jv�Ü��
i���hٟ��i����<��^�����s���J��]�l����tE���{��)�eG��i����1��`��I��(��Wv���>��Z�v
�HA�Œ�hS��Aȧ���4`e���;_��_Z3S�C�d�Ξ��m������0�.�����#�f(|{M ��T�Z�Q��{�/uȌ��I�!uy)쀬�B�|G^�9�E�r��!�!����N�� =�v��=� k=��f1 ~�*��5ioksKv��GH������|N^ԙ�Ǌ�`X�� Ai�O]d2~t���4$8�%ga��v��i�R	J-�+���q�s���"���u�u2��C��Q~�GC��5J ^�tF�3�W�VF{P
�3.:%�=_p�g�bj�6r�ܬ$�pN��F��B}r�>)��?L�n�Q� ��p|"=�2���E� ��Q6�	ɳ��M��|��o!�*���Ѥk��9���qJ�iK�!����ʼJ�	e�癛��u�$�P<��������
jg�Ƀm�q�hcƨ-�tHS�l�?��5$��\ȱZ����gؼp�"�oԓ�_����(���j-[��°'Q�[h⭡�u���@�҅(�/�̤��$�ѐ�8��j�������Hh�Ը��%��:c�Y��|p]ѳ"4��t�/9�Ȳ�L~U�`l?�§M=ى���=.�nɊ�x�~~S�A�)��	)�L��3���^�i_�ZO��wl����!%�n��=��x��fy쾵K=6�C�J�C���_2�h��p�Tx@.(���G�V�{���9}�m=�!���7vAN��	�"]�4���C/�-��VF-v�]���o���YD����|ބ_P��]��/}�=#���9�:�� Z�h	*�ĕ\�$�Y�zH ��։/8=�H�a#2쾆HV'����u�胶g]���̍�xI�!z��Kڻ�uB�q���h|>��"���<2T����a>-��.�?��=��S��T^�ۇ����]j�w���ť�(�Ԯ�3sD��S�>�x�F�.��h{g��f^r@!\^vgp�'�0U^��și1���j���nI�*�߮�1�к:G�'�3��cB��N\i�`
ŭ=����P��!���pg[ ���N�@�\.��h9DGSn�M,%����D\;�
'&r�/�x���L���^ȕ#��^ˈ�O�kz���\�d�P�_�pT)^[�
Uz��'�D!����Ј����9ROV��ݢ���~��{ٟ��آ*p�xϩ ��c
3�/�4�A*��wAk4�W,=�����<�!��`2J*��!�@�b�
�Ə?/e3�! ��Ͷn3���[WS�<!>�0E�2#�!-XH��~tD�
���mޢ��f��O�v�l��<�d�i#�jM�	e�X�rL�#�X ih-q�;C��6��m9
�S���״T�y�:���βu��%��W�c�����`F"˸���c4z&:vƧ��m/�\������i�Q��o?s�_Q�P���V�9g����eG��/���r���{/揭��w�Y�l�9NM2g��ymǘ�[c#�ё7�oDG�X]�H�"��s�Y�	���T���Dev�q��Ϛ�Ɣ�
2���I H�����X]�`��rp9��?�)[���"u�R������v��R�_�"M K6&|�{]�Q�Ԁ�iP���d3�����
Ъ���G�:ѲL��i���v΀���c\�8@�@�������S흒�-���M��}�h�@�P��Lsǉ��@�Ƨ/�l�M���	�hj�ܹ���:vfW��{A���c���'��T�Q6��*��@x��������=��>Q)jDc9Ʒ�[-���x�c�S\�k]T��>���$.��(Z�q���s4-Ɔ���Y�r���x B�%r��!�S:�?k�
��-0�c�O�&����� ���O����&Hy%.��,:m��J�xCW���x�០}in8ȃ��	��@�$@�՛���[�����:&���;D�?�n��P�� �k{0 �|;Ϭ�q٧�0.0���='��?�w\O~��;�@d��6�Rd���!���lH!�m��9n�Ĕ�%_�qH$2�ᇆ�<�L����m����G�\�(�9m.�Ml<rRMt�˽��{����8�Kjg�4�vB�µ��9��Z��g��w�ƕ-G��)�v�A]WQ<�6R#8B��]=u̓�G@����e=C7�/3� �ė�s����
��9!;�K73sQ�h���f��s���8K�Z��ݻw�8T 7_�6	�ѐAâ���w�!{5��z�	�n��2Ch��.`�0DY�ה����HS�j�-`���8�ܲI ����������xT�J��54,���[���HcI�Sr�A�+_���-�	iXK�ڠ�a?�گͩx�8����m�u�k�g֎���c�w�d�-g�e�w+�	ly������
׼ ��A���A�"IJ��;��>QU��2q��qS���J�u�@�|��D^�F0��f��HuJ����>s���9'Ba~zq�������"�3�b�e;x&!%lk���\��ۏ���YZ'�����7 `��(����w�wG���6�]�#4y����-���_УV�U���p+L��@D�1��d��tWs"���JU�.�l�����h���ϟ:}����-8ܒ:g'�����$ݜ8�興w8S	CW�f�FL�r7z�&����晗OX�sb�o_�ۮRy���� �	�pEEeeT/iMtS�+�q�����c|}�sU��m�����(H�\�[��M�]d�5����b�5�]����+Z.w<�S�M�2�(�*N�1�����h��P'��������M��ȑD��E{
m(�#�o���i^'狎��ks|��h��|hrmC{���o�������I����nx	���ݹ�v%��ճj��{��o���&����3K��x�R��0/��qe:��v�PD��A�|8��{�ft3���lr�щ��!n��J�w)}}}J�nJ��}�R�9��#�@�{p�]n��T��5ϛMB*~�M�|��ZY���u/��߲�_�Z�^sIh��JeC���o� v �pM���5�
�c����z'��~ym�׋�+�@@��/CG�b³U�%b7w0���C���\�)Е�|��&��k�e�*�m-xx�]ځ����3�n����t� �u��K�*����� �}��o� �¾��\Y�yK|	�z+��z����r���=8��j��N m]c����R��V���d���'p�s	2���6��H��9_����Ge%�&1��k����P*T´G ����vn��n�9��;���?@�Z��ܪ���T�Ӯɣ�d�(`9O�J�X��W��9�rǪN=r���Y70�5�+Zx�O/mN[���#��.����8�v��}ϵ)ٷVf�Ǡ�s}�H��f��F��a�@�Id��Ӡ�����G����C���D�U���Є�B�D@!��QX.}�Б�¶Z�m~PK�W���B����d����'�0`��T��w��\"�������&�y#�i2�������c�*�Y8*s�V��㕿�jRl̳$�����D��S�SU�Gk��)�.�ۄJ���`�9����zA��G8��� �G&�$b��9�w#�r�׏ʚI���9zB���:Z��2��~L`�(�D�>�Ԫ��_/K#@^i�"�#��
�&��6��{�	*���H=��I��R�kbЍ�y�)�84򏟻m�⅄�ap꪿�,"�/��M�-��
��O��� �*H���0 J��:�7@�"rr����7�/pOv:�
m`&�&�c�pa�I��mG��x���ԉ�p���
���5_֮��t��9�� I��6��7o>�@p�NM���`�zd<�߶@�T{\Z���XHP�%��u�7�]�9ҟWƝ��Z_�,y�ie�\]�}���m!zPe=�/������m�W�����t�-:a�G^���0{;�5��W��1˂^tޟq_���wlA��{#�F[V�ҹ-N)dGF*Ȩ(L���}^�	�����3���W`bj@+6�^��,�xx�S�x�;��l�:�v�L��@�Z�dǧg�>�T��_�í�tw��?3�GD�*�,p^|\U~^ }��h5���	z�PR����ɳ��d�+�.	3��{��A$�-t)�_;H ��h)����*������ԍ�?G���;hai�0��*O�L��\n�0v��۷�x� ��˹rg�s��/�ޭ��+��A���)����`�t%H�怪�o�oF���G�Ңg�$%%UӨ������U��x�%;�P�}ݱ��'��9�y7�6D�n@U�A��>(��uߤ�/
S�WF2|��?}���l�����Հ�7K72��(��w��Bt�/���8�a�ϴ�W<��Q����n��� ٢�S� z�%�ː*
�������?����6���\r�V5u��A!��� :��PR����G��X)k���tM=�I�$'�c�yИ��]�KB��|�]��5B��m�m��*���5�b�m�|��Æ��+ڍG,h��M���r�O��RY�Zh�M�@��,��G����~'��a�F��Ի������
GB�jEq�#��*-�T��Wo�l�2c)��ro��g��|ǚ����W$�����J��9Bc�E��ָ �X�X�x�Ω����TV�~hM��MN����'�B<�Ğ���I�%��"�d���|A�C{kO@,�T�3PYJ�ڷ'/`0�	�w��M��-�׿#��Pt9i"w|g�����}��H/b�g�i��]E��!��z�W��Ya9�5�{�e�.vqaT��`ٳީ�b��y	�y3���;8�C[�}̩���@�[�vP�]*�)Rf�a���RnM7c�����k`�Gt����e��h�L4�["�z��'��n�; [UlE��q:{AL����>�B彶���Lmk|��ym�ď迊�7���������e�!��=`?1֠�� m��$;��BZ�h�g7�����ĭ�EAe�n���+���
&�y��իj|��(	��b�5��B{�g^�i�n�(���smD�qvno|����KC*�M�gcc�6~�4��I}ڌ���KlP&d�1C��
��;�/����4�-�U�t�t�Kp��:�%��zs�b"�w�`6����_P'}v�w��ڠ=#j(�)N�&�S8�����*�C;���r�پI℣i��'��h��:��.��i��˞�Z�3+����>��==
�R�F��O}���E��ND�*Zڠ}5��-�ͧ@s<�%�U�E&{ OBHѽc|MJ�I�i��m|:=C�<8v^��P2���m�o��n�mv��&�<����,Օ��סʃH�!R���~+F��{�^�Յ�i��
�D2S��N�A�7���xx��;�m^��'��d't�BєqPS��:�3 �s$���1^�j<�Q�	3����E��+�D�bҩ��Ԧ��\;}����M ��'��?���v5U{^�W�`pd��/�ŏ��n4YgŢX�xV��%��h��채2sy��g�>���7�N�S��=�ro_��k��4�v9yO�uvr
������9o�:#3�*IM����9�]�C���C~rwt9�d�'�钠��Y�K7�_f)L~����ۤ���w�Bͮ9Ƕ��Q��	z��c�OU\�yU}{,K��5C�v�������i��ڑW�%;gƮ�H_�q�Gqh5��ؓ��p1'u�C�~�^MLT��!�+?T,o��?v�����5���C�e4�e��=3#?��=��6Xix6/[;g�WH�$R&ZSߏN�D��+^��;�3���u���e�'���`&�m���oB5Qh�D�jr[�����'��W\���&��h��m�5�wzx�c�^��F~MӘqzk�z�9�,~ґg���G�9|_c�[Ԡ��+D+O�D~��[6+�qS��M��FJ��X�؍�C�YrK�#T�UL�
�M�u��΁��hC�Nۈ�����3�@H�������wɜ�,�[���a��M�b<�܀�H��p��o������({�+��B������mbpk}���!��$�GE�2Ԉ�,~��k�E�Sd��W###6x{UQbf~~>��u~1/U#��0 ������r��o2!X
!R�z���	���j��?��C8���*��0s�M]4�;�/�BU�2��ߠ���)e���S�y<���Dj��L�g�Q9�ӟQ��vi�q�*O{W�>�`*r���q�I���u6�Zę*��u��z�ם9/9�4�l�E+�)/<i�{&6����������(g�����-�6� T�5=8j��D ]����{i���f��Gb[�����c��I��	��SOC46�D�i,4*j�Z���^�������Hk��L(��"��ڔ^�	�ƺ;���m�M��������R�q8ףm��N0Ζ����@�L���\�xAV�j��*>�r���/SX	Uo�8�$\��@f�q�oB�t1�K�s":z�J��}�R/K�{�RU6쐈/.iS!�?U��pD�T��XV׻����F�(�R��O�|{�r�����n,i__��jT
_�}�hZ�A�&�Pg3��V�
!x���ՉCFRw����<}��̖\�1�����8�/f���<���)�D.�X�R!2�aɭ-@ޫ�nd�����JT$1t�^�l]�]$�C�
Z�LN`wB;��2;Y�޺� }�P���d��j}$ґs@�{fW��T�N{��S	��� �S_��+i�js�!�M����*��m���޳��dj6$�np�;=,�<���}7�@W9�vĩJ�罄�1�{���7���&x�yԘ�7*꽺�?�4~��W���B��$���7o�,����@��|��[��c�g��~�~CK�v��l�w�j(G�$LWzvr#���)���E��x�MH��n��zC�4���G�iي^ǂd��O��d7�j��"�e���h�f��j�B�m��!�K�U��;#�#a'�j�*�0��ȯ��׳��(I�p��mM����lՂ������0_0�t��PZN�8�a%�_�
r���j�8�7�?緜WKpy���S�"�If���i���S�S�ހx6R*�;<��5U�z��tq������h]�)I��9�Ӱ]8�e�e�M��M��eO�^A��>�:�[=+�d<Zop�p�P������SN��.>�M�������*qA]t{�ɹ�$���:�N@د�`���{K��#ϲ�t�s^�F���%}Gu'{�X@'��c�{dV��'h�cd�&Fٳ�%�I������L��gBKZ�����ai؟�}�+;�?��dz_�Y+�j�[H��M`��\�S�U���vѩ�H�c�)��k�A{��h��S�C��z�Z���hf�T	␭�`u�$�D��ˡ�m�hL����-�����W���[kP^��(�����=�����v{�/Q�����yhM[ܭ2�S�zw�y^x{��vT���ÞR^�TG�3�'}w�a1��>: �N�f��s8S3���NɵlAG�(�f�C���HxZ�2R��ц�����;:H߭�E_9�{X��H���Po�GE.�����#(�"�^���ŶO�z��/��9���u�.�Y��yV0��bj5m�4y�n��&9�����;WT囷�D�7��B1�����s���k�Ӕ�"Ϥ��uʋNU��k� ��1����;3���D<�`:�[�7K������C�E������	��6���W���;j"�1��Jp��
�UT��!4)|��?����_��D��D��ֲ�7�fe>oL�Voϓ����GiJ�=nCv��y��ф���Ԩ��W,=;�������EM
�{s����S� RG�{U�{RU����U�V����I؛��w����N�� '��;�x��3�v-�C6�ɕd>#�s�lL�''`.�]����t���w�q��E���Y���b�m#<��֭R��Y�o�l�q<.�]4�o��w��Cќ�������I Kk�ǃ����qܣDZp����n�ᚭ[�ą��m����n�C_塟�ۑdі.��*��dv�6�r��c�j�rt_�z���W�}�2dꡫ�=Ws�Jp�BWd�Ѥ.��3�ɔ[^ ����h��mnX�K� ����D�
W6��es�:�yz��k]n!�� �q�N�<�0�i��8T�ǘ�'r��@1	q�a������3RhFVS���s��׸��n��=�����2�C�(]����mZ��~�c�A#z�vptt�#*���߇��m4�_�QS&誦� ��-�p*�#�˟��K�kh^i9d���r?B8=*6����$9�յ�z ��&�I����Օ��˱#�<�I��O�k
���rձ��;��Ӟ�)�NY����C����K(����ڠ�Gb�ϑq�U��8|0à=�R�,���=�!�Y�M�XtJ(�h�X���h�^�$ONJϥ�c?�����<��O,�є���`[��?�<��� F�vl�&4E��p�y���Э�-2����%��k�L��"�ſ?�-ɜ�&r�?���M8��M�A�n$���7ԧ�:��z[vS;�\Y����׬^
=P@���,�>��L�X&�_�Z��Tu���W�3��}2Õ="7��]jzX�v�	M�(|o�O,
x>��L���aƔ�H���
�ė�\�;��W9���O�]��Cl�=�5�� ����}l:�+]]]	~� WW�%�3\�AS�"B����݆x4��=�#��0������%}�G4�����C��
���&'������o�OԱ���h���r#�U�@>��h�����(�y��� k�^a� ]�ӟ�~��˰����Q�^!�����0@ލ<��o0v��$���4
f�0���d����fM}��8��n,�)�ŧU���� lt��y�3~�頀7��9i�c?�2����Bȴ�7�H�#eO!��"��"IZѠ�2�_�&W���7o���3��x&4���Hcdu���� ��G�߿OV:u��!R�!�bChd�Oi��|��	lL�#?�XuMP�O؂��|>o���=�s~�%x�+'u)�:�$l�o4{xxT�`����{����24�w8���|�K�2�G?;��	8���nN�������^�|AHӿ|���l"jz�K��"��W��@����O�ɜ"����Y{m9�3J��&9~x�"SD�h���1~1��2��4�����U_H=�$��/���/��3j*�3��*7��4�J�.�|/��K��.��7<���z���~RuU����K�v0ޢbִ'i9�rf��g�.����A������m�8�=�(�!y�!���hᎼ��=fs@�*;��.�U��fS��~y(&�<N�I�ܴՓ8�>�f�Rb�%hn!n�A4�wE�&z lEcĸ��w���@��H��`a��W�n��0�C�$	��5�~��C�'�ji�}�v�xIa
)�'ZvgDՁ�&w��B����æv�x ʝ�٢�c��6�O8vN�b�0��A>���|��3�",��mE+�UO}{�J��Ҥ(���{<��@9rR��L)Z��q�L�H\�����*l�_`�V̵K�+m�f�e���h����ÌM��J�GR�w}��\ׁ4��1��W��C1D�pV>���p��=��:���T��(N�5"�D�}��Xxl3�4��ox��j'{��?��ag�����sT�����n7{����k�M0-J9*���l^Z��_��}�˗�'o�%J�Ю(��cSI���
��6�h� ]��{ܗ�&�~|���:��;ft�9Ry���/�5J�E������VM|�$v���S��@1f'BW���T�k�G��͞���K�P�� �Z$B����ۣ^	��uD�sKT��}����t��DS\��t��8�2�W�&�2&|����9�|�:{�Z\O�LLJ�1G�Q�s�\���G��'�j!n�(Q�,�$�<#�y��E�B�RW�DH���>.;L� �p0+x���\-D¹Â���9��b���6u-�#l�Q;q�����G㶚�Ł`�'2jԶ��
��,H�T�9��/\r�dEL~U,�R��Aѡ�7��%r8��u��D�&�-���ы��#� ��t�3�d�%��{��a�Uh�(��8A.7i��v�)xޫ�7@бԈP�lo����8h)E�%�mW�g�+;��th�x�]-J���Uj9{T����P�q����/t����t3����&vj]7y+_�=0�R�s~	h ?�؛܀KQ���G�Ll��|������/�.�{I�@�ܳy��uاȀ؀�6��}�ҵ�����
H�(n���{�����ע&��j\�j����$�~��|}�=�rp!��@OS�p�@���2̅:�e%���%��B�������nD�k�,=]@���}�i=L��-���� �;�����wH�����Fo�t�736�ʱ/��MLG�.�=��r���s�(�߼qꔑWK�l_�f4cn�#�e���k�����h�ɗ�t�w�5%xFxM����j�����&Z!��AX�tA�`˛�1q���^�X9�/��i��U���Ǎi���3�/$�6Z&�<#+k�Ͳ�ծ���=:�6���+h����;>�v�L�!�S����Κ�(wlr�z����E�G���{�ծ�y+;0A���g��><��&	�(���H/��J�F�$#Q�&cպ�Ca���1�:�2}���>��V��o�n�=u��O�6} ���>>>3�����f�,�`���"�B;�;~^�J��M$-~�~w���=�����9��\����Y�}!����8s�%�h����q}����(�6XM�mMie%�n{����r�M�щX^a�(�6L�n0�/}D�!�)���8e�Gn��#	�l�{\%Ϗ�� s}�j?�m$U�t��c�ܩ_ �^�L��y(�p}l���nz�R�iU����HK��ڋ�C9Ż�0��E�q���Τ�%�h}~���Y�:0֊���X5l.F�G� �s���=1	����91�L������44��D{��'T����Z��^���`<JQ�+a�!��Ρ#�L�`���d�]$��&G�<%	��FMM���Ĩ���l D�75���nBkt�:B��'����0�>�;ohhz�'x��d鯩=F�����]g�K5�x�^�ul�ϣi�9�*Љ���W�Z�ć7���nu(fب����W��X�l�����P���}g��.y�\�Җ�C��zn�T��ccc����2�|T;4���C_��'CB�νV��3T*������|�����=f������jK��B��hZ�n�ki�.�ѡ�mgFބ��T���LӦ��)��_��s��r�n�ЀΡ��C멝zy�=��Ao�����lg��N]F�g������R[�[�:�?-/<��{`��i9�R1��A�<������0I���V\�:i�R��T�"F����g�'x��6�g��o������ڗs3#^{  p��+/�h�8>�h��a֞Pb�.Ȫ3Ҟ�X�q��-~�"{;x�L����[F��kuN�^��Z�M8�fה�OB&�������t��z�:_r���_�����3���S����
Y��;M:EK)����S�Mm�^;�~[���.�nE�0T��0��mO���ݘ�b��.��/�%䦣2���w0b��������?�o��H�K�jy%K�Τ�k�'ԳF��`D`��g"��B)3��ee�34����jMiv��W7����h�(�PZN,�ptd2)�(�+�nv���X����=Z�߱v�
pf&8�qP��o#F��$6�Y]�Z��}��}��I[��+��xn)��hC��9e��kߧ��U�0�t_;��f���h9x\�k\��|Q�>}�Pp�f<rF���.BQP�J�\��d���Ka�]-J% ��T��2يk@�\�,2��Q�_������A1��g��D)�*�yC��/�	i�wV�$��4g��p���ݟր뉶 �𧦕ձ�U;!HR�]L	Y���}m������3-�����wO<��n�i��jW՚����}�
���$kDQ��^�J�<J����K[ƣ��z�u2!�w�q*f��߇��KZ��Q�P�	�ড়P1� OF�L�u�NL�}�����Ʋ�5��Q*�~�dz^�f�q�{F�<�3�[����B ��r�C#r5�o�^	�g����!�dx��-��PL݅�>}4�x z|��M~�X�$Z��� D���b3xHZ<^���ŜߝX�LvP0�ۢ�у����|��v�s] >-�P�Nk�5g�­kK�����~�#}X��q�ͮ��>��[�%g3�4=������{���5Ԙ.���
��������Z�:�,�O@��q�'��ح�y��I�:Ѓ�z�.2�l6�����I��[d�-��&� ��j��Z]1��Sy�p�ƕ�;a�[�q�ѤL������<�5��~ק�GM�8mn���_�l&��-����_H /�����L�����k�)ʘ�߫���z�SyWHT���q�C��X&q�}��uk��J��ϕ�~K�A�PL-��lWd^ý]on��8�T.��~d���1�(�(d�S�&Ɋz��c/��W�<틈aQס7� �-F��m	$�͗R��$>���Ӓz�^��K�xe��W�W9��_S��Y�`��3��|���㹖ȖD�� Gt���QV�: ���R�P���=��:��)
}�<����ѡ�o�_k'&&lJ����i<k=�n%�D�6��l�Y5����+���s�BA2:��z��W���Y���*.�utC_f�?��
�~�)��P%�K���pV����=��"'�EVw�x�v��}j� �Gvy�t�o[c���,���Tn�⢀&U��Z]Q�rސBV��W�,���)ˀ!�c��2���01��'�($�I^�����R)A��@*\َ{CE����7 �+�{�7ܕ�(+~>�jG�υ�'<Xum�f+PE�-���^�΄쟸A�p��3Q/��}�������S^��Ρ���ה��k�Z��0�Ïo�Ү��s
_�����*B��Z�4���3�,.Љ�,��%��o���������sI�̔Bg�*̤��yڷ��U��� >�*Z\a\3k�?����V硿�oE�������M8���K�^��#�¥�]��v�`�:���m��Ya��휣�b�R^�i]wD���Y(-1��h"d�{m����5k�U�������Hw"'��7�`<��z������D�O������~>.����#�ﴞ�_�'�����!���F`۬�]1*�)(WIY-+B��2�rL/� ��c>�N�`��&��e\b!	�����ߥ�6�(�l\�v�tq��/���5���xe�*j��)�����p�^���Hs@L-ߐd��C�����
k�'m��]�[Y�^0VO�e@ *]~ ��5���"�	���)��j���Z-Pve$r��"c��Q��v����ޑg���)c~���p��|z�H��Y>|V�K>>nG�v�t�P��Q�T^�2�۶����
�1�/T C���f,��b�� Ib�Cq�Q�7��^�,�K��Z����if� 竳�FqX��S�*Z�,����c����҆<xSO�p>,grz���w?(܀H�
e�����[��|�["${����!r�Άƀv�be�W �-���������3gu$��/�j1`u��q��?����bE2�P� �f���Id��B):��N ����+�}�
k�6��f����v5>�靁H��@˫�9�P	���(�XB�Z!���[�jXJ<�]��`�Ѡ)�v���l,F��I�)��| ��@W�1j>c~���ys'��i��'�M6�9����?!0�C$�8E���D�(��a]X ;p���"�3�__m��`��3.]zO��£iJ#�^�C����΋��=�[���AyX��?+Zě��74��*���4�:�[G%�s�y���M��|��(�m�j�� aԞ=�4�0���r;�3��<��X�`TZ������L��m��@�{5Z^���Rؗ)�ԏ�l�ދgO�O�t��lE�y=��U2;y)�4���^5.^�%��,�G'&� �ٯ�Y8�s���/{�E(lp, �������F�뽇{
ʱ�s�㹅{�+�S�ˆ$��B(0����]�����|wr��,��~�v�=�'A���y�,���}����0�n�|�u��+�D�u���çQ*g!�Af?"}���)E8!$�W#����e;�T<ic���>�O+�N�uEX��F@��\�Z�E�4�ߌp���!��ЏӦ����9AO����(����8����/ �&������Kjg~�(�Mgo��R&�WҰ^��^m���S`�:�f�{|:ς@�-�{�.�D`�?�� �mF�������aB	z����Y1[��lG%�r�D��Z��0�@��:�[���[���M���:B��\n�7�l�N�i�}4���3�H��!��������߀�tm/�k|��Њv3䡜>/x���|U��A!f#��ku]��jas�F���������0Y�9�xZӁ���-�q_Ѫݑ��適>�ղ���l�#����O᎟d=��O=����i����y��B�>�ĪO��?�������<Uσ;�T	ݻ�+fg����mL4�@4��I���L� �3�d���
���2�#g���?a�Ⱦ_e�9���V�54��Q;yG��/j"�H�ajg+�՗�@�C�k�V�nuZ�f���_0����f7��4S�E��$�1q��e,��#�1�r�n�S]VV������I��`��O�Eu�:j�%�F.<�C}x�Զ���	s�r�5�oA����Q\�%��6Bh���wA-��l��� �8!�g$	�&��d�����X+�+����>S�xd@���\E~�Q������̡�#9R��}��������}�F?�NϞ	_�6�|EtȻG����[*fȸ�Z��J�l�+1�:-	��u��0�gB�hFT�@���kh��1{��Ay�7�(�'��Jz�������ձvLL�`�xTr�#}��|oMħ�zy�3Hu�O[�@SH=n��rq�E��m���Z^�2L�O��i8���zm��~M��Ѧk�D�/\��"���ˊ�A\��'��:��P�l
s�� '�^�n@�\9�>y�=p�+c�����r�cͼ���>b�Cp�mA�?���W��B"�J���>�5�p	����ȿR||��_��5�]�Fs��hÉ���A�!�RY�l����N���7	Mm2.������|��0K^��Ð`>�1.� �.�~�a�Zi�-��2���x{mJn�*�束�O��H_l� ���'A���E�v0���3W@�נ�׃!<t.�垺{b��ub.�W����ne��&�A��K	�9ϐi�$_U�C��c�� |2�\���Q�H�0�g�ΚC�J i5�DW���#�q�xᳲ�� ���zv=>Nh��c��ߕ�����j�4?�������-i-�I����d.�����Tc�dVa�w1~�=�9�:8��1=vM�l���(��x��1kroHA��p�#��mt��F�g���U�w	Ew�Yn�U�!����>j'h��r='롸N��mvlI�����k���:���Qu�å����d���{޶I����s��'�����S{����F?瞅���S�(=�bTV��.]A=I��n����YzV����|���2n�:�ѼQ�Y�&�#{UR*H�S�q������U<���-��@��-{ݬ"���v>y��fX(np��<���W�N�ko�CWK+-�E7F�H�ӂP�����+�[X1Ÿ��kd%�����SΨ��d�#WO~(��EΝ�?Z�oٌp�t�T#8�`3{�0�J�����d`Hq![=�<��r�!�+��W]�)eS-��;z�<��,TҼ,~���Ktg ��ڳ�o�+��J�Y]]��`�v?��*@��pU����ޟ�S�����4h$�Q�J%
E�ШdHi3��%)�$TN���쎐�:Bbۆb2O��Y�Y�:�߿���^�w��~����p߯�u��{����%��K�o��}ς���PͅKKP߇�b�XC�Jh,�J��a'M�S)��k7���J:�|�f&�O[��h����
�Do`E�%�Ⱥr"���y�u�ڮ�i�L���řV\K��H�E�dIC��4�1ִrW�Ps����9aM����{%�Y�]D��ޕMu�jY�[q�Խ ��]�;�m)�F��!�/�
��j#q#ٺ���Q��y�vXta��)���f]&#���É`�8�M__!�.ӌlxB�'o���\�ՖEtdІ5��N��ʝ�'���=�],v�tw���Hl�K*��t�ZD9���t�0�#(ԓ���ͦ�1��H�:� T��t���:���,OgJ�h�#�1��V%ئ�
�]+H!3/�������Gtb�:$t����ŘH�6���gf�4A��٦s�m`���R��:Y�]�ҧ_9gpVk���\-q�?�81����������#���w�%�C8�FS�PA�2Q�ѓ����R�k����&Ժ�LS�B����v��#؃͋�A$���1Ã�:��9_��^�g��k��<?_��I�Θ9x i�.�Y���+�9@g��Ϡ�x�(��3��$�&�v$>y@�I�!�e�fG�ڮV�%��IlN����W��O�C�Ğ'���?`h�Ǔ��z}+v�=�]��i��Zsf����[E�_�����b����3��
�Z�x�X�y��a�-Oi��jc�f�}m�tU�0�2���)��T�X�`1�v�s@Q�(:���XD|��@g/��y�j��"ZF0����/��C����G%��_�?dr~�$v�r1ֺ�a����&@�����`YR��ŏ��%��ʣ�=�6 2 zBm-NΆa#���H�e��,B]���W�g���I
'���.��'�b�Dg�k��e�/(*���ق�����8�Qq�V��ںM��)�,η����\v�����ӳS�.�������'d�X��+DP?ڸ<�jw^�,��S�>�A��c���i4�%�y�F��#��3a��	8�)lSU`m�3.(�,S1X�4���U[}���.�7y�>�̾�_���5��:��j���4dp ���Do5�[d�2F�c�"1�Vq�j�cdb�ٸ��
J�E¿�z���3�׍�3�z�1i0��]p�U2��q��H~S�B�B�w�G�"�
��*�{�?f��h#�������	���m8t
������M��0,xj^�<�e�#Rǯ��R*�qV��4B���]�[��l�:x�ʻ�Y�Q��y{�L�2�}��X�u�v�	���}'P�������@I=ϿɈL���O���Y
�(�<����M��C[�T�z�Lߊ���`��H�����DL�#�FFze�H�
�2���@Q�7���B�Io��!J�X��b��Iڴ��ӹ�Q/iS>Q�_�0��=Bh��i(�Pi��T+��#�i��~~~��*_����cۨ�w� �)9?�G��e(O���Rw�&:���=!���=qd<,�zx�2e�xł�2'O(�^�!׊��Ǔ楞��:� V������j���E��O�Ǒ��H��]�&�T���V������)���X�Q9J��-���ߝ���h'E��Wgo�J%� Ü�����y����%����8#�$��viT����y+!����rG��VA��I�E$��n��n�.�S;�&����Y*�x������ۙ��'���kb']��-t�J�
��~�%���7�˝�;��o4���Ź2՟�W��ؗ�L�����XG�|Mw�^w6oq(wP�K����(h�/_vOs������f����ʇOt<�y��l��t���ӵ�S�/+2ӧp��7+�/w1�z�/lMc�����}Ip���'� Ǫ�wH�5���>J|�蓶���5�Yo��㐡��t3�\��ʽRMK.�ǂ	e�m^�_}�7!�Us!Π�o�ܹ�f�f�P�:�f!����cT=P>��u([C:e����o:�2��;`U,�υ�+�^�ki�2��2���A���]�m�Apr;��>gǊ��+���ΰa؆��7������m�uO��������_HP��c��>�v��R`�o��l�C�����cLdz3Ф6r�8՝��-|.)����KX!ո0]����E�7N��-��=ޝ���P-�Kq�<����;+,�$b����ҁ�錓HE+ksH�������w��fd��$��˕'�?�ܫC�|S,���CNx�y���N�Ng)9��K�Kc���o�瀧���.�?�3լ��'��u����+����JNE�#A�x?##C����=�(�ؗ���w�~S��E�t�K}}=i.�?����c��1�� �GCV�e���_�������@��=E�(�m��/��h
�.�R�JZ6�	9̆�iCgg�OۂC+�B|}ۖ3����V�����X���1t�be�h���R���	%�ju��� ^t����`���ӵ^������9�.�Q����Yfn�&j�݇T��j�H{V���TL,�Q-M=�!s5�C-�����ɔ��<B�c�I�)�g'g$��1���o���k��	J]��<�l(9���C����6\���	�-l�z���>^��9�ӊM�/��%�=��lxD:����ṛ���կ,W�k�P�]�~���ٽ�=n�ߪ8��j���˛�w���\!U���Ef���2̚v�yυV1�[f�drQ����yv��u���̯��?w%�)��+�;����]���]���j�ΣL��Xyl���������i��xC0�\�]�]��&(��F>���x;0����qΏ��狘Umtx��`|�����Vg�@�B��y�)��ܼ�,�L���W�hP�Ӓ�?����s�Sا�� Ã���\�˝oFz�)(W�ǐ�-%�ۮ.'�}ؒ��_lE�$��=��|Y��*��oM�o/�`��+M��\'�'�w�W�@>�qt����ѽ�Qظ]N��a�=[�6���xԼ���>����P�X�0�5曆����v�w%1ӵ�{|�m�h+��o5!�_K��P)Ͱ�9��9�n� ���WY���pִ������YC���R���%ў����o6gM�L!����T�Pp[�����o������k�G#� l��:�j����n'�C����2���� �ڌ������8'f�L�Ȝ�f�r������{<F�r}�L��7�4���x�����9!��� #���BE(�ր�����辅��~ju@�%`�j�풙d|m���d�lS>���#s�m�fΥo���M93\�'ݍ���n�Si�֮/�%�&џ����Hִ����!oB�y���Q�zJxq5DvcP۴C��9ūq��7�t�>J�_����(����8H�ڸ�S�>y��H���������t�b��bF5Ѷf�R{�4v�_�K+��P|$Z�m�;ў>�f�]_8����X�f�1�IK�y2��}�>��*]�«��-�	W��:-`�M�Hv��F!��HS�&b�8%&Q�̪��[�pS�v�o6�l�\��ʜ�v����N�������C���BA��Y��#v��SY��⼇>�}pZqY�Q8�8��j��BKc)S�A��@��^�����]0�O��s��;���]�QNv�ei��)ĈY��ZϚan�꧓|�.՗�J�:wLĲ��	ɢ�?�q
z�"�[0��]��1g¢r�k�/0P ���4�fF��M���I:��WGQ�Yf�{ �mC�𯴡&A�CXE����GCv�.,&R4�<�1e�tљ��e�2������u>FN�	��WG/�a��򇶢����>^�>��y����`M�TmqP̊�n�W�q������?�1��;��v�	,L�~d�.sJ��(E ����5u�EQ�fY���i��:�`}\��T4C�c#���v��w����Œ�J�p�!(�q�c���Y!����Lm��e� "��$I$UXm�d���&$�@	�K�����c�<j��W�>��̌%�5�J��	 ���ӟ"e7��ƒ�;qХ4YԱ�㥯�P�@ˊ��)&�ksϱA�A�r�K��"�������@b��>F �O�����~3�)��9�`���ǗL�9��y�{�A2ω����~> ���k��m�
ʘ �m���BL��;�.šXsoddĂ@w �b����?�:=�ZeV|{�)���]K[.!��_���"܉}S	�B��`��*�G�X6�h%�����G(dv�y��N����9���u2�ξ)���=�6'�_P�	B39�׆��1����<�R����g���'�pS�
�;S^���[�+w���K'm}7��"&l�Ӽ��A�R�N� �v�X;u�l��֧(�#{�^,��5;�Q4��l�-$��x�sw��������]�>^�y����,��$�(O��9�ƿ��=F�K��Y%Sf�C3������$��e�{�W{8��im�}�p	���V/|�KK�ɓi��]qj�L�5���.#�5���|$%&s�=��C�1� ����Z~%�2O��+��$c�Z��i����s;�*�,�	B��rR[������KBii6۸4��8��)It[�(�4�F�;��&�5b�kh#M�3��(���wn�>lZW��?:D,X`�"�H#z:�|\���{S5�Ub����b;�����\]I5͝�װqF;e
�8Zg���X_�@��6;��HEWC�<2�(:������~�ߙ�KO�����yyy��"47�$���������0��[��[��Ry�h���F��
E��;�f�>����@�x�2���S�^�XJ '��`!�d�Sʚ�� ��ϋ6<��uo��)��J����u����6�K�o��-��%�����K>�$��}.�����o��-��%�߿d]Χ��d��8�k�,شtQ�k	�w��'?�9���NP����l��b��/�G���8�E�b��դO]���YS����I3�a������N��l��_��=w�=����_�����Ԅ��<�x�΢G�9�X�x���xYeŻ�p���lʷ��Lr�W���'��+�cC3Uߥu3� ��X��%⋞k�r0m���F����+�
�/o�Qx���H����=�0����Ig��I��Օ(D���u�'����3̓��ȋ�&o��}7uss�����L�n�1���ϒxmК�N�:l��������L�M��͇$Ѓm��.%��1~�;��Ï�S�u/�X9�<��kj'���5�r-�G�q�o�+**X��sx'N\O�u���fr�����|�����!�x���߾~}��X;���e����	�h�Փ��O<w�ɝ���>������!��XK���&�`����yy'���S�=_
�ք�������'��3�6�T�VR���/�?WH}nP���G�w�
�M�7|`ZC���hu����)\+#q��;�sVV[�f�]mt�'�����c��]�����KľL�q����޾w���n5��8�u���())��}l���>�����<��%�t&O���Ŗ��$��Dٽ+��s�c
��z۸F�]+�g	�0�����ݓ5�L�z2w��Sh�ME�*�՗s'����Z���m>��K�~���4U%��d�](E'�<����Ν����Y@��e�zI�K&����`�/x��X%��ܖxhZ�&/#����G���@�}_G�����/gg�E��1�8�v聘�ĜOn�x5U��[kIݲسg���7K���{�ʪ�P�j �h���ۄx��U�yRNJ��|֫�3rK˼���HI��K��+6OP
*��W���}IYY�>�٢;M�:�}�$��1�U��F@�͍����1#���l{�
�]���RZ �=�j�٪��u��a�����x����.��'$$�$���i3�6��"�����ay�w�=�<�#��t��|����P��P��5�p���YƑ/⍿��P�T��L"W��^�H�h��}�����¢d�]�=��t�Ѹr��"u-��K�
���N�
�	�]�FX����z�t:f�0�3yx�Ҽ��ɵ�����������W
��S2k\�򭶬�Mc�QV��t�o�uN�Hԇ�"��5	��ș qCR�����Ż�Yj�l�c֬Ys+�Ħ��� �`9�$�G^�g�2�Y�y}ʑ�	,� Iu8��j�+ٙ�����;�(��}��á�D���,z�֚彽�1�!����ew�0?|�p���=d��5�j�[Z���;1P�rQQ����_��"�R��h>�'�ؓ����g��QZVV������� Y�,�Nۯ��C�����E��x4�^�xx�9Ȅ�܉����x����v)H�7 O���d_y A�	5gq]��V�%T�-n�U v8�i��ݻw
�`�����H?	���e�4������ڊ�F�U�gj;;;���y������,�r�'D�ꙃ	N*�$I�l�䜳�@���TwVXX��E�~g �/�P�=f���C�s��ȓ�ʩ������ɰ��k��ҹ�o5����K��8�@���Y��\>����v�)l.�6ـ� ��l$"a�H�����>8!^�q�"�2���ֹ����꠨�"��و0���6�����[�D��kп�������UZ0e�jEp��Pҫ�4�*�77���;�(�����_o������&3D ���_�x�K��no�N����>H�J���)������V[FH:u�C����g�G^nt�����_�ǲ@Ą(��9�HBy���c�Zw�\i���颦I�y�!)���l�o�o)�eOw O��׸�e�p]�V�U'F�}����`u�h��j#h�8aE��\��I��
9A����~�@4�u��ȠT�AX<�a�?}}}e���5i(�ӭD
�Ҋ�XND��F��g�\q�;��?u�#Ȟ_ӧT�^��F�D�/O,vPШIZ�0$��XG:B��s���ψ���G�������\�Ȭ���Z�S8Jڎ�6
OĔ��p�3���3簦�8�����`_�l�$�����K=��K��Y����zezhl��� ^DP糳�S��?��z|>��
�����+㇓kX��<�Y@���T��c�����	3�F�ӹ�\�����dw?͇��SrEݜ�?)������X��X�|#��8 .H��.z���ϟ>�vR�%t�p�51�c�%�������s0���'���NЯ���Ќ	�Z����_�F[
O�6�a����0o����(i@n��H��Z�o	z9-6+s�/4S�U���l&(9���!�-_JN<���%H�6��
��Z��Ʒ�ՈWx08��Z�=�����	�����ju0����~��[|IFٖ��������|�>b����?%�>e	.�qV���>��V��Rɾ��Pv��̿�P�$� ��{&P<�d2&R��ƙ�!�(h�M7>"�=l��F�;�NG�1�"#�4+O������=_A��Z��KI��F��0z�\r)��V�t�^<ovtt|x�j��ϗ�9c/�:�Iݸ0�&-H\��SI<����j��ӳ�=]]\��IjD߲�]_�(��-�l�PeY�_����3�a-Mf��|(`��� ��<�{b��5
�q�[�)�9���<��]X$��HpǕ��ֺy�~!sI@A���_�&h_bz>D"C\C�za�����P�BfZF��cFF�6�#��8~i%?��}~����BHpH\k���˗焊'B "<�㡥�l2����u=z.��W����B0"W^k�����߲�ju=BGuʈ�|�߬A< �?P<�3���2]P�z+[�����U�m;���o�&:V�	e]�_[	�J���u�\,�E[ֳ2��4S�ѭ�����͑���D�e�SI^y�
Ƒ�e>h%��ڬ�0J�c�Z�٫x���0�[Éߕ�:q8�7��
�: ����ε3@?6-�hu��"�����X��y�p|����=�`��f�sX _�G���sQܐ�3ӎ\��O���5�m�v�@1�����7h��a'lE��`����Y4=h�C���	�$��P���Ȁ�%LTM"{��v�#��R��i�lBO���S���nd����c��pҘ�U��ЎL�M%g�h���� Z��v s~�\ �K�Q�O@ �m����J��@�/�<�qߴ�w�\n�Q�AS���|�o� �@����3}�RG@蜟�t �PCÉR%�A���N��p��Zm����D~P��x��6�0�X����$L����P߉��kyAb��SS����$$?w���E��-m�D ����ƴ8�Լ6�p/mQ9�b;��S� ­�ʪ�<��%��,eS�<���+��\4�301�<���f�!F�Ӏ��|��K;ہ��������G�Y�ś+a̡���'��$�SVvp8�l�� ��fNc?+##Î�7tP�1�pI�M����8��|X�q7��p�f8s��������1ϒ��o ��^^^Q � (ـ�,(���\%��m8z{��K�){{{;gg����b�yN�x��#vt,��U�|�! �K'�}�&�P'Z�PE1p�t*����u-GLjz����ȴz�'���T~��~���Qd ���|T��\N�-�̾Π%>�.k�d���5B�p%�A�b���<Fm�LiZ���\���5'�[�Ò�eAAA{F}x�S��C2�(-�$K�s����x��1	�7������gTy��
�4��F|��Y#��8`�����	�Y �g���sEX�j ����X��USR�K��Z�3��@q�z}P?ꛠ
e����e��_5�����j���L>�&�/P���[s�.�1捞6�w����ETDd"b��H�p[#
��䱱����p[,�@heq��+9g�8�UI�;Q��`pĆ�y���hsf����nNN���C�M��p�7>^�� �Ċ[Ʈ +;���L`Ts��MM�
�\�)��>yG�T�t�)�g�p��_��^K�t޸��y�>�tC�'x���֞#)%�IƝ����?Y9d����@��m��x�u8��V���Y��f6���ڞ�\"XsJ����%XM�f�!BΌ����?`l�Wu���(k5Z���'p�ף�f�&��!dw��[WX�BLG>�_r3���-?:D��!=�PE�e��w��������=���}۷����"�1�_~ �DSq&Y���:VHܴ�8��&t�F�y��g�-~d�%>��ضe��%��P�YXX����1=��?z
�)` ����BjY�tYY���hޣ�,�f�'�I,C� EFH�tΨ]FR�,/�b�D����͓��������3O�bWW/�
N}I�Kh�@q^b�&b)S������\mVP���Q��C���R��,/����]ڰ�����d��k��Czu��@PN2��8<KQ{�k:�O���0gB����|*\�/9��28��1n��MT�G�L�^� QU:�WUH�d@M>m���"͎���/��ֲ�xВ�ɏ8�GQd��gl�l�M���6O�t$7(B$)�?�VX<��_�I*q�'O�o.	+��&�Eo���q���#VA]Э{� 1=*��7���tz[��W-/y�% 吺H��#\�'Z=�<}]�f/R�)ݍᤴ]�.�1MnO%�8�+���9V�a}Z.6�k�__�H8��gh��Юh�#�:(�Qp�[�,��V�At[ �������}�
Tx%���豦��ka ���"V�5�^�SO0�J���9IV(��r���Ff;�<��K6:�&ЋU_�F���t>J
 wW��w�R��y3Pdځ�h5R�ǝqrrzO�l�4b�jM��.��[g�*"�"E�T�֊@��X�j9�N�q��2��Zq�j�	!wb
�c� m������<��K���p[&��j�� �yJ�r_���	����a�c\�P���#w�(#��8!iZ-��8���G���5>�Yپ_t��ĸ��xv�����Pe���Z��ə2�Q&�����[�?����{x�}�4�b��A+��C=h�C��`w(½���c�PW�����eQ���i��k�3�S�1���SS?Q�v�0!��oUD�2��yyy�'��o aXS��܃�e���4���Y�A�o�6���6���Ci'���;�##�j&�BB�c�;::��������^�)�-�ide�_ī�q�����6@��$K (�Q9߿U%eDEE����S'���M����42[���@���W.�����>2`ooo8�D��Z�/Xs�eJu~G�q]'䖖��s���x^~~~&��<����VWWǐ���(��	�[W�e���ͳ��/����8J=ej�/�A Pt%U����a��x�����J��$:��vǓ4�+��(a���S�œy�'z�	&9��� `�#ěڈg�!�Y���8	�!!!7�S@3��pg��	��ё`"@�&�~y��w��PHyrJ6���r��ǜ��B�ĨD�)){(<�6L��R����M-�Pϲ:�:,���b��U/�rw����ꉊ��Kӣ��'�j�~%"<(Z@:#�<L�.��#e�l�"n���h�9��[`,�Yl�ᘱ+C�w�v��c�qU�ZS/�a�I�s�.��?�k�iϞ��h��p�S��p�r�3��3��3><��F7Q���y�����.���!ƭ��_� �>�$w(C�B:�viA��Lv��rd)��������B��&����Ԡ�FQ���Tdd$���@�����X,���*a(�R$_���ܰ*y��4t��	����H>�r�Jf���mkKX^LLL���F��Jj��� ����	a�e8q�L�np�]g�?��`��.�o�}||0�1S�Sj=�t��8*! 	͉ll8�p]��L���|�O�ƃ�\��"������)D�IS�V��Q�>�ycw*΢���l+
��޽k���1#��J&Ҥd�1�'Nl��	B=����b�<�?�`u26>�Y�m�܅�x�:���<�	>�|�\龸p�_.��}vt��_�����/�Y�����}i���+^|8�W���T��{�$2<<gC��8�t�НOt�@�V8d�>�����[�Ŕ��^���?��p�9U
�[ww�a<���ד�Iii��N�H�w�*+QJQ��fy�'T&����f�l��f�A�6KrÆ���ʄh�Ș]L���29���"��f[AE��왭H�����$�u�)�2 6�>��{	6���%ǌ���-��(,$)�P3���144D�*�P��l�'�рqU���fnnNOy�2]K�!(����^�����e�C���'FRa%͖�2��Z��g��@{a`��šq��]���ߠ.Ȓ�T�݋'��ت�����o��}J�N�X�c`$�ܥ���
tk�H@������X�q��o$ZgS7���[F}P�Ћ�n�@�l����
�4�y:�]I	�ܓ���ʪ�	dޥ=�!�yU��u6��POS�hUU��E�%��~w�����v��b��u��l�0)��������Ap�^j[�/x^��<�Adt�X����y�v�eFHH�+����i�e�}� �Y�ٍ���;���*����("� � �
<���@!�.E8ST
g(����h����^YY��`0DvGiwrJ��|<*�s�ܘ���`��*咖���Rge�m���xg-�e=?�^*VR�p-c��ى�X��,���A	��0���̰���qn7J�S(�~Qeq�H ��@L�0����[�B��kEd��������* �����MފA���a8���;
�vy�`�VBBB�Zu�����zks�y
b��
��;)�q]�T���ɭ��t4�P���0�ɭK�:
[��$G���rѓ�[����B
=���(_���s�b��R���&3�(r_��h�A��o�⢿����Le
P&���5VVVw�\�}�H�c~/��u(�|VXX�	�&���@ſr�d��&M�UW#�@���"(	}���5���Ζ�~�/���dan���[�&��$�Y�%���=��f�T{��u}�� �Q�SX�S3NWRp����2Ț��3���G�[�D=i��z����75���T��F ��:��w���85㢂n��g�_h�ۏ��m�4��#��F�u�>J�&�x6d� �-���QY��Y����?��/?�`��|�-�"�iuP\�elMA@#��y�������&���/�ߓ��E�=��<��]���j&�ZB�GB���p^OO�~DO �/%%%ɓs�0;/���M e{SX�cF/b����ւ��B�Y*"**�Is�ޔй)����ၫ�s���6T�3~b�� n��_�G��N],Ėc�9��!іd�V@���>}�l�2u-��S�+���져�|�L!�����)�r�{zJe�x�;�7�<�Ig.�^Sb��␄8���F��q���h�ԭ������k�95� �S�11��Ȃ�@�k����LϿ��z�-]��MK���/�!$��������FAK�A-9eC���N��s�\��x�[j�s��A��{�6�� KB(N�SI̤�^p�'�?DS{{;V/�H*"�@�JC6u�?�6*I�9.��]Z��<kj�2j���͛'�a���F����,��o:f�p���\�
J���&M�uc}�<���R�-)i�8H��AW�A:�:�����Ɍt�*(ෞ����~|�J >:��6��ņ�ed���܉Ȋ�+yu��*C-�/C��?L�j͔��{	����r�^ ��k(7�4��$V=�	�U��ng��x�@qܤc�;���_�*�jkU��*jĐ������&L!�� )]��$+�E�?������p>�_]�p�����d���hˏ�]��㸮`��"u�����It��
���i��y8���f{�={���7$)���� 1Rx;B�6T[E�?Խ����STYY��8��i���kvv��^8��n��0X1��[�註�ɓ��H�ߒ6i.jř|6��5G�ʳ7/�OB��)�vv��ĩ���Y6�Kq������kɝ���p{944�:>>��q
�,Ζ4}�=cF��l���c��2Nx�������)������c%h���J�tj:Xt���^�s���� �3���>cFRYC��EM�hsNk~o=�M��RK�����"꨻:q�Zhd�_D�$vU�vu��
�-����dƜ�9��ܩ`c|g�P����:ܱ�����v݌2��@�(�;�R�[���}E;e���BB�ׯ�lE�!P���H2t���+�f�+��4*��胢�r�AH��������
s\��#,2kٲe-Ǖ����d�C��-	�v��t�רm���(	Md:T���čj����:w��T"��>n�JK-na�T��fM<�X��%,�V� ����iOi!�ˍ
�0����-B	d\�3��LF����1��G�\��eu`%����B�����.�P�M��8KV	]L�t�vnAa~����F��� �(��ʧn#䍠�,�~(R�=���fc��������"&�e��*��䯽T:�|l�+�*}98�h,z��Fc�*��E�;J~$N���[ϑ�-���f$u+,2�c�Us�m������P�Z~&y;�H������>��d	��ɘ��I�,C�QUPQ1DwlS�.S�����W[m��t�����I�f���Ѝ�j4fs�����86�v��딅E���F��`Km>|�ø�ĸ�A��u����d��Ý��;���b H���%]I�~`�)��,newi�Һ�e���~.Vl�NQG��� �R���n�����a'���DP���PE���� �&漁�???�-^T(>�#�uQ����;af�9�F����J��0&�:�!`~](�Ѹ;�Z,�e�>��m4�Z�`@:,3ĉ�j����P���� ���
��0Fe�??�I��j�o�����.��r��-,?����i���Q�n���|��.
rT���u�0�y����$h��ʔ�]��X����`��S�U��pm�S�P�� �hHS� �(�ni>���ゃa!���mSb���8�oKS���V��h�|��g�I-��dS�YJ-�������|F�����W����}q�f��uA`�S �A�������=�+9�2��`���F�F�����}H���H�ڈ���[Z>N���\��X!tQ3����ͱ��/씱
g\�-?�]RR�0�9�f�P���n� /��o�@9�~jRC-���0��F�E��F��<�e)Yp}��3NǺ�x�������f�jx��m��F���N��l֨����@{
JJn�p2�>�AB���#���b\�a���Z�b�Y���N�]�J��j�Lvs�]���W8��')��;-�s�]�~������ҌWb3��7t��y�A���r).��Z�mgt���$@�CЏ��{�pRL���!(555�������
�E��'�_��t���(�ۻwo����_H`��dd���h�q�f4���`��2gv��r`n?�Nof�s�љ�ϫ@G �W��N}�1ണ�cjr2�G\�ǣ��3���J����c�ݨ����JR�JY�7"ԸC?�ΏE)�9.�����\�����G�������e,5G���~*�M��CU� �
_gq^��E:)���w�Jbu�bG������ Nd�}�*��P.��>�4x�d"/��.�A1��F�V����W2~*#�E�E'G}H��<h�f�����d�k���erB��w�z�3e����e�{����}������p3�L���XRJ�WWYT�4w��|/�.����c�GL8t��h';� f//���˾rT���<qpwA�7r�����g��,��۱�����H�rRr��\=��0�1?�@L�����o�g5G����o�z��n͓��P ��W�but�Y9KT"K[<������S��#��������v�������>P,�� �78������s4�eTʍ�_m���,�_9G6t_΃���#��s �wU'z;2Rt��Hڛ��%$��֔3q�3���k��mB�}�l$B����K$���&��� �nnn�x��n�OhM���p�g��+W��%W�b�{r*G�#��S1{���[��w�U�┉���Q�эS�d���	0����?����P���H���G���P�&'�����Y46�?���,���.f��S1�@�����IM�y2T��b���@Y06�}R��ɓm1B��q9F���#�;�er�9�a����w˪݇CӘ
��C��1�l�N<;-�i��U��%���`����^^#sdM� �B Ta�s�����IU߂���<5o55I	�s���/��֠�F|�\��G��w�Śs(u���1%�I�'�F����	�(ऱ���`�J��P�Yvu�;|���	C+u͕5%߾Y��~i�@�!��# �L'�i��=������G��3Ô�jao�U>���S{���s.u��Mʺ�~�3Ф#��
���ohhPp�)-8�8���b���MT���ԥ����@������(��kMv��;枃��� ����a�Z��5�2�Y�zU��޼�Vi��P�37�[#e����9���L[�#�d�ɐ��S�ټ;���Y�c�����n2�"�� |�N����":RJ��p�Z�����_<{�i6k��ʷMv�R��8�8i b瞢Yk�x��
�b������Lf�=����,�_�?� d��k30�t����DmIKo��ĕ@#)����minc�㋠��N��P[H"�')Jk���L�	�bpP嫑p��1�oі�ѭ��wO��ߌ	C����������u�WJ؎���+u偑��Ē,vN�6\o��N5">����T������w6g�D~��Uw�טn�-���l��$Q�BX����.��(��luhv͊�oy
���Lg[a"�@�
�F�eg]�=�������1SH�Dtrtt�̃!�٪�*����-��E�����g6�N����\Y�#�g�:�!�RF����!�lLLLSY����m�;��"/o�u����������6������!PM�����H��<wvvVXF�kn�N�e��#����iH#���
Q���Q�ub2�:�
���3gC��a琒���ɭ��c���n���Q��bo`��m6��7�5Y�2,�N�
*H<��ġ[[��	O5l%6F+��}��U�N\�5�9K
����,��A�Ȯo
5D��x��0����k[�3�5@�q��\A�T���c�;P\}oP8 şξ�2#4%���(b�&�d�^'�P��i�L��
m?ť����-a%�iFH�?�� ��[�1�K��y����<�*,4t�G��N3��X]]]�@�Z�qR\������O�*_��n�ƞ���]��3��
]���ݨ�1�RI]��d��?}�*-)y�␻!0��3�N�U2�c#����Z�s	&9!׮]���	�C����s��ul�*���ɬ*�-��8����u˚��ZXvǾ:(�s����<1q��O��.gZZ�e���7�(~T~�qwԇ�sO�n���p<�>���(���q:�^c���ju�|n�FP�J��/���f<o*J�˶J����8:9�*|��BI�k�-1�p��0�Z�U��"Q#U�wGݠ�Z�ӈ~�m|x��*mL~�LG\��d���01.H��O�F�s[���~��VosW����i��|(���)�^�`��]�I�|x�]���szhx8����vŤ,�|w	mN�P����#p1�ݎ⪟v;�9νh�>|(���S�f�.q���zFF�>��F��H�&�r��O0S�� ���?}Z����۶m�ɰ����Ay�����f+�b��I��t�d)5:�� j���HQ��7� P0r�j��ǳ1Ϗb�׽*?�l��+d=ř2QlNA�:C����IV���qɞ?����)�?G_*�2]��<)�>�T��"�����U8[Ҽr��&�~S�a�w���u*pa�sNYD)���@�N�8�`啼�]��;g�-���^o�o��J rA|��K=P(0�U[���K�ۊ8�(S���'~�8%7\n�}��Y���R�0cU�ћ ǀq���ޭ�o�b=P[Gg�)��z���iiU	(W-���
i*�)��*����肂���U4�riiitC�xdVF�9ɽ��2+>7(�ڟu�c���]:uo6��x�ړ}c��o
6ų�[l�ɼ�|�w#�O7�/N\���xl8�|��ݛ��8������2�w���B�+V�)�M_�h���d/t_�(~������/_�|���;��x�L�;IjLl#���,}���;���MsR�tx:T��cN㥆�4��!>��}9d�c��)4?CΫtp_�n�JK�v��ƪ۶�k�%�U�.l��cF�3���vySs�/������nm�B�ۍ�eѝ�sr�V�}D������P�S�c�;G�ٜ���.o��~}�a$5fJnl:��ľ�z���W��]��۷:����Aj��j�W�����"y�ګg�B��i�9(�G���;����
a|{��!����o�������w�÷���u&����Zf9l��K��:7Z����[k��>�\ڄ1݅��ͷ��ހ�_�y'�}r�s����d��&2��@e�M��99���~5��ֽ}>6��oP��.5�	#��
���>�,�qv��<� ��3�U4��_fd��{[K�q]%�l`|��q��xX2��PoKR��,d�s&FF�I�S��m�@����aٹ��*����v��7�p�4'�=�|*b��cVR���Z���c�߾=	�9�A�@Z�,
�55߽{���uF	��ú_�\{������\{h����Ȉ���䋠ht�)�u�_3z=sTSr�����8���KS�g�svK����t��܀������!f��Qf ���y{_���ŋ��7\R���:�h8�|�ңŤ��<6�)<V�A�j�:e�r�	��~��e�aO�}$q�n��K��e]���#�ء�)�d�>D��D�G����IS �i��v'����a�z�PZ��QIA?�T��Ҡ%��w77�F�� 7�<������J�𲉿�a����`��d.��I&��K-�CG��d�M���N�={6fS����.�?���-If,��b������3��[-Q�$�Ӯ"l�KY�Cv�YY�J �_��j�"/��"��2�c��q	��wa���V��\��2	2L��6^���,&Iu��/������R�,N�O6b�ݦ�(���B�w���@��\l�J��f���Gƞ�.�����F1r���w�ܴx~�ڭޜc��taQQ'
��>��]㿀���@�-��O�Υ�����mD��V��o���S��c�B�̊�CSU�%%�$ �3rK��\�e����ߤ�Q3.�3jk>�60���%����}�;�ī�.DBo;�R�� �]RUq�rµ�ĩ��9��j����A�O]��'��J����0^�����2�2�+MvK@@8)�_�o�+!C�ގ�ᶸ�ޖR�HGo�-}�Tx��27���b/SRT'�rr�a�sw�Y⿛�8�4~Ǣ�oUI���ሓ����9��§�5�2�X �q�@���|FqW���(�yvuu�"{u��؛U��So��!��FJu� ��c�`��ħ�x���%/��0�܍��<x�`5�KC��杕[�Ғ�	{���������u��x�!_~�Ҏ+�4��U�sqI�k�P�$�3�CK ����}A�:��ó\?����գ*�+ �Nɬ�5�4coj{����|����8��CME����y0��A�JI���s�'�d��HI^^��#2wx�&;#A��zkC����2:R��]�I�|�ͨ��
��9}h�=aTϽ�7ⴃ��S�晑T��·1GpHt���1�m�>��[���G9��n�[e�<�� �q[�$�b%�d�޽���G���6�<H⤤8-:Y�m�Ɵ���&����q=�3J�SY�\���^���,�W
������I���
�	��\r�D���j�Ԍ��m�y��%$$�as��3:im�*�� <B2555姰=דz�������}�d�A|$0�c����~���e�ov�b��A�P8��4У~�(��2V-}���U��4�����'��*D�wp	�	 #Z�`�A��J����:�Pj����8ݠ���R�ۥ-d?�n�����nn#�E���a������p�ӄ?��}��m9UI�JJJeX(��X��ء&�ii[�Y��/8WX�ϝn9�W�\\}3��:{(zjrm�/S��ñedd��1�H���H�����TfM'Y�&f2}uu%C�[Fa$ �����N[��K�9�� '�(`6֟#�`�el���k�C$��5����dK��7��<�4@*�nR�v�^�����,�:����sa��j�-	�.��7ߎ���Ɣ�C�ݴ�K�X�!����	{��/�(�2�F�M�';7�S�&���26�7X�'��Jnnn��Ҵ̨�SD�	��訨���(�"i�Y���QE�k�=��ɺ��bbأ����(qY[[�'���d�j�vO&3�4��������b�!�8�b82DI�I�����S�֑���m�NF8�sv:+?m�u�L7z{�����0���D�$��pz�%Tj8!�)��ۓjg�υ���k�Ki))nz�D?����zl]<���M�	�XNS�R���d(�B�_��^wش��L�M�;$�����'r�{�p�ǀ���?cR�'�*��<�K%ۺ��[�(y�@���t��0��<גl����5'�����w�H�_cc#]?$-/{/[Q[[;L�)PwW 7�viW��Y��[i⵭��gT��:�A��/o�O�H�UA����	I?E������P���GZT´Q��V���(��W�Ț]F�'KSI�[�ƒ�����aJ��
�G��ނ~���9�����/�}����<���,�s�����̍���L��p��4�z����v��_�	Q��۫����_���� ;�{�s]J"��[+pwj�@\Q����x��ͷ��x��D���+o�ǿ���[.x��(�yak�1{O����(5־{`��1^���*�w`�ث��B*n��S+�w����$�OَʀΊ�I�-��������OlVB͉'w���ɚ���G/�2�����7G�#b�� ��g7�|N	(o�f#|B�x�dS5�lq�"��l���^"�ߒ}���G׭[���߭�b=y�u?� �4W(�O�nĳ�_ޯE�ree�E3�#k�M��d[��x�/�0��<`�4�^pkkkJZZ�	�BEQ��PR:�M�v�?z�A_W26𗯸�k�XK��O�>���=Y�q���(7�X���9�.�Q�NB�9E轛{"��Ӱ���\Ł>Cu;�㨑d�/��8�n)�0�U�W&Q(�F<�d�nR�$�
nfs��4����M���]]��� 4<��7��0PR+A�D�Q`�P.���Z2n�a�6^^^9����a�#����^�"����ߛs��3l����ب5ۼ�_�!���y�ga� � �~�b��4^��]%f��Ñv�n^�PD��.Ĝ���/J�����rq��c��Q�jR>I��A�+�mn	{z<�b��~d�b���X��]������ؽXzV������z�� d/�]��&�!����5�p�s�zn��U����'6�B�@�|�)h����p���+Zt���aX�nb�lsWD���-"��R���v�qb�V� ��v�?%;(���e�l��rA��Zy^ ���Cw��bܨ2	�f��f�"�~��Ͷ��)��+�I���{�����aL�Pn�O�6�s<(�Kł��kp�f�����v�oOyd[IP;��l�=۵1�M�¶u3��(	3.o=)t�#>��< �S�T�y��k���d�u&S�%�qHd/�n}������0�\�������瑧��*�e�B�.!�b��ح��?{^�5�T�����ͻb�y� }��É�Y؆��7���ěA�O�1��lq#B=��u�u����؅�3�=�Z���PUK4�]{�ڶm�7E�Q�r�XX��]x7`	e��G�5���5~+�e�
)l��^g�g"zI�Ph*�� ȟo�Z&(��p,�y���-h�孕3�psN����W4h������Ӎ.�Q�|�q#�3�>�X����"4=���<#(`D�������I��\��f<Oj�	E}�M��2	�5QUchV�-�VB�2G��ٚ5��~붉���~iI*�������`m�al�bD�-B���)w@f5Z�<�s)re�Xd�����V^�t/Gbב2�CO��7�F��6w���z^��
X8�*CU��CQ�z�A�]��>5!����铃W��F��"�~pJF�r$���ʾ�r�-Z��[v#�	��5=����
�=C��ODZᰤ��T�ķO�V��l��"�d+A_NBOV|��9�1c��{��En�=l�`j�g�A�/�rs���+�x	�^�GL��=x4Y ���/~RD[�эj�;�Q�ȝx&a�s?� ��D^�{%������� j���{L�<<bjU:��N��"{��M��������In`�cUUUx����^[[���H��ߔ�F�}$x%�{d؅˴���pD_��(�y�˯_�ЍS+� -���qy/
C�H�[��63�mnn��k�F��y�D�P_n;jR-�'��
� �ݸ;�yH�c�E#S�L�/<4��o1'��<y�2Q��C@
���M��0A��M6����F*"z|(��0X�p�r;b��8�yب�]�ty���M��
ٌz�G]H:��<>�H�&l�sIlZ�,��J��sm�q�,��7�ܪ�Y~�cj���`�{?�$���iy�,7�+~A!�0*%�e.6O��z��tLsGu��ː���Ti|���>�9}����rS�O.�l6)/����[�+ ��}�8m�]��xIA�K}��]�F�D�������(��h�'ZͫFPs|�"H>�Z�X���q�8Y>uC������C���(h�K�i�㘺��+���l?r;�>�P��$���+����;���]��������E%���]1|�}�T%�)ytd�l���/��C&t�&\.%�WM%�9׽@�ElS`���䖍>l�`��8l.$���ͩg���bc���Ԓ=Ӫ���G��`��-1(��T;:kh�M�� mT�i$�ȶ"�uu���&괪��l�x(co�d`��bȍ�Z�����|��`�?''��S�.c�4�\��1V��o�C��|�;s	e��IQY�x�����{� ��;���*��m�հ�sswI����f�C�[�9���+$�ʮ�V�ݺAA�0�q˘����,ǚt뢓߷"z}��ωcM{2z<*�ܭy����ȃ.��crjMTi���	O�v.�Gl�z��.���Z �w�WB�0�Kt���mgV�A�VF5ц���2	t<l�oA��Fnk:Wz��4[�o��F=D�͋�j.��a�=�ͥ��^W �s=��)z����!Yf�x>K:X>���D܎���P-}V��M�nz�J��eۅ����-AGQ'��Q��;g��o�v�Z ����ڸ�ǈk`�m�eQ��9�8e
w�)���^�F|�
��7s j__.�,�p�w'�����/i1D�I���̴���A(k�:��$�މ�D�Jx�sNl:���l���q�<tw��fQQ��Ρ�HT���=�sY���U�=f1���-���i�^��f���K�zNd�ǎ����62J����w���λ?$��Z[[�U��$#?����bS+H��?��3y� �d��d�qww���5�ޡ�-��2��@���#�5*Y�-~+�&ê(����phc�Ygo�>���B�Y�����5�(6١�
!@���x�Q���6��ˇ��ՉoI�u�w�ō��d�=�*v{$��B��h`� �1G���~Xo�_�˹�J��)���$�з^m6���`�]�ws�U��`�Q��\׍C���+sh��t��W���4Aa	����}�3@Y�~���zJ��4m���z<���)S��^ے}j>�Sa��YA>�s�ώ���R*��`���_�~����#��ΐcT0�"_籐����Hn�*���늖hH_Q��T��>z"�s��-S!!��QZ��4����������]B��Ԥ������3���=�-�������	b���á�
D�	�������@�Y� �5طg�Ac��f�U��x8�n�y��j%hFY�+ƞ�y8>0}kLOa3�P-��LP#S�3�8�;�*UR������)�rP���;� F�w�3���y2"�3��WG\�y3�����@y�P;ޕ��Xt�7&m�������N��"�a�}�C!��s��Bz�V��ړkQ?����1Q���OsA!�d3
_��*�&�ay+�V�@j�q�w9��E�.\�
X��/i�g�\ga~��c!�_�_�[�Ե%��������|�/E��)�[\u�1O�!k|�=�gI�����w�G�V6��555E�YQ�ZW:���qcwH���[_Ծt�v�"D���|�u6���?���N��!�"
����EW���A�}�{э	{���<R��th�� C�g`q0�6�I���&��h$~X(��7xi��}j����uttl���{f�ֲ�j�������$ԧ&��B	�I	�/�֓�>T;�a����ﴥ��jk�98?9Mi���	���{����5�}ſ<���8�m>���gyܲ(X��B�i	{Y/�!f��ϲ5G��wT�j�cE��=�n7Bf���[�94�����%,zt� �u�c����ϟ��v�X�����l�t0���誮��O�IAq��s����DeQҘ/}���h�(1�h��g���\�աR
@�:�DMd�o�@|���ؚ���3s
��\#��j`u�͏�6O~~���dSK�/w�\Ɉ^K����Yk���_�G���n�r��Pֽ��}f:#�<-�kW�(g�呁v�vH� �D���J�H��UE��u�5�M�����$ ��d4���$�c���$T�µ��k��7�t{�',��X>��Bs�A<�nY�������IJO'52C?+�C�i������v�/���t4���n%C��q�	֟K�c�褭<v��$�� ���(�݃���/.��)���zg^18ZQ��=�S#'����Z�4�s���k��$I��{Lq��8�C��z*�h_ߖ<��5�{<��]�*�؅/�sL3��,z��WJ��gc%OZ]א��&��"���\"��w�d1�PF��4�ou��	�������P �ʇx3��i�V�w-B�����.!�U#b��(������6QN�~�¹���Ѡ�V�� [�Ѿ�zw��k!�X�$��b��N�PaL��쉢��;�{Pz�r ��>��;lb�e�v	IC��~sL������OtjN���<�T�7:����浕�NCA~c�~Mь�?{�o�l�ӘAEC
�;��J�<��y�0����V��X;��_��}�2$8�`{��8q2����w���L��7��
Qhc%�]GB�is$��W>\��� ���R����ѫH��-:"<�`��%���+�m��r���C�M6��^�0ٚW��ϔI�F��Y�g%쏨�L���d��وi��5&��v_h����O�]��d|Muu:f�GҪ�א������Ʒo�y�N�"9���|�� �lR��ss`�����K=-Q���Y�:g�_woٽ�Tp�����+
�!����3b	m��:)��~fc`�`��'K���Bm{woQ��W\i�Ȋ���[��ͽ&ʥ:�����6��W�����4��;��e�ꛑ�}>%
A"/��uaL]�\Nm�*߼5����7o,���J�G�S"Y�����Ʌ1��2���z�C�E��\�iڸ�AUB�R�WP��=vS(�O�ݢ�5��� `����R��xr�����+�-g��<�&����c�h�[��Ѿ����g�
��X��p�:�+��v`D����
�S�ACeeecG�\<f�lQ��'�\���	R�{��+��oT��ن+�6�S�_W��w�/	?xv���􈶪�Y*<6�.O}�0��cA�f�R�_�M�J� ��9}�xw�������F���)��M��-@��4ukM�yd�H�w}o��p��[�����r�����w��6���,}=U��j�s;m���00������o1��
��M��aN�(�ns������Evo��^�*`����~++�����G"#�	c^$g�4|�P�^�W����V���!��n{_�c�]|8h8K&A"�T�	�1T&n����Qϊ��ʗI0%���k�RL��G��R������� �Z����nm�,w�a�3Ӌ��*�/���r�9���&�gL����&�tx�ܸ<��e�����<��2i(A�q�Q�D�衙�YײXm�sk>Vǩ�&W����q��Jl]E�o:���;~R�H�IE�Z�B`�6��J,�+���P}:όG�BcZ:�<r-̇(sY{P<DMvN�"E�R5�+��XE�����E����=ܻB?�t�U��0�p�`�h�h+w��.S�OG��ey9�뾚���<߁���~�
�!s,����(D�l"�=��Zg��=���
���G�3p��?@Ku����Rj���=_����^����L�8��k��^��i��/�Hw��(98я�G�t��
�|@�w��X@����s\�s�2/8R!QΨz��r��*	$ް�lM��ޚX����mn�c�Ѥ�O[��n��|ི���L=)p�����Z�-ᝣ7�~�:p��]��:��B����&�W}�;;]��R�Ie�xc�&�"��f*���lח�K"��[�U�C�t��{\��g�MGF�t��I��Z&�¥�|
[K�Ъ��x���K	9><���괟���P�d��y�����7*`
o��!ڷ�z̠P\�'�*�n�(�q���U*d��2���V�$��`c��3;�Wƞ���>f��z�p��n�b�E�j�O~��!��d��y�GW����}�St?-�j���u��_��̑���1�2I>����^ϓ>��*�J���]��d"���[��W�V?Z�Q>v~�Ґ��澚z��aa���>�
�:;��������Z[�k3����T;C'g��GcY�\E���1tsd�{	Ꝕe<�a��4+��e�|��-l�~�c�E����9(/�ۦYSZ��D��TE����X,�&�k,]�%>h��G��e���S�*1U5z���HcX�6P�u�v���T��]aU�q�4�,�-l���|�0��^־�7��~zW��{��ٍ.m��<�>�X>ͣ�j'k�*D���aG+�-u���&>��8�Gs���=�bt{k�4-��խ}����������B�x�c\
��9�iU�4��H�n���@]�=�N�h�5ED�����T��.�B��Nf[B�_^�kFPy��V�G������G�m������X'�Fcxa�}́�"�9�̺�Ci���(������s�Ѿ_���e,K�;�t�	�|% ��c�ij�*�cYn�n��*��\6��Y�k�UOKɤe58Ǘ����pVVV��W-"��#:21�{�v�dk�j���HgK"f�_��	��̶�����Vd��Zt���C�PA��1�|n���cc�49�\�kc!n� �i��K��b_�zf:��%D����iT���,�χ,���LB)��|J��<�pH�r\�	����8,�����x��H��Y�#!����A���g�L0ݩ;�.w�ws%b��6�����Bz<@O�H$	�c��yHp�]���hk��ЧbW�qow!��:�'r#�S�����p7�Myw4�1]ey1����j�鉪�K�i�FM#����i���=��8,i5�%�����kac�ϊ�h� ����ސ*1��_� �s�b���4M�Y��s���9�����ZK-o���P y�C��B	e{$�r����Q�'�E��l%n���8"��X�bUaв��[)�1��#亃��J8��d�P�J�S62w+������6V#��v\3r���ۅA�+R�.Yn/U���飏Wz�¸�o�%� ƹŬ�e^�]&���=��EV�
��i�j�c�$ �t�n�>�+X��ȿ� ׇ��,ӌ�	.Ó�G�0��J��!6t@�o@���A_��P�QOXE$kk�%ƒ��I�>���J.�MoszW�I!����:
d��m�v�r��$�a#6U�^L��y~q��xGEE���;��H�K{�1?{71�Cl���t�3p���T�.0_o��8&/�K?9������Ǉ��Ch�m�R�T���	���f_���lꝖ"���Ȏ�J��l�=�P$��-�����]�^��)��K5Q��8��w|x܄�R(�߸�@NJ�*���.I5��C�����o 5����k�Bs��H�=:2���	�:?���$���l���*F�D�&ʴ`���ÎR�c��<D� �-��[n��o��0��"p�_��1aaa֩�[�G�e��"S���u�
����+v?���}cIv]�V��["��U����ׁ%�d	
��A0m��Ph˾����i	�=m�����'�s�p�~@/b��)}U�� ����K��&K���*'i�q�.ʠ	 %n����������gʺ1B���{��U��L���^ z�ZeWd	�b{��`8�³W�l�Nt���?()C.��c����Jqs��+�}Q(��bbs8`jB��|g��P(��3n�r�A]T�)���$�I��".��"�|ZJ�s��]���E:�O�і�tT�Q�t�gx��.�Î�6��1�i���m�;����q�X�$��sQ�p�`���OGF��s�([�	�:7�ֈ�~] ��ĥ���v�����⟜�[C�Z4���X�/�T�J�+|0�޸[���Įԅ1!���Uօ�A)ѭB��EjXt֩�����-�W�g?�У�Ix��=EW�^u+����c?�%X��xB���IbQ����{�*�fi�fK#���GGG����X��WB�~WA��W�:��&ƜU��
@4����?Do�%���i������ɡ����.ז=�s�NT�
$?�L���n������w>��pOF��J1Ns��nb���9q�PfK�r*�aǋ*ҩV�#ցPt!UX\�SRbt��3���3�M$�L�n��
X10�����Ę���#� ڣ7��q�O��z#��߼R�[���<�T����5~�뚙6ڊ^�	����.h��z�VT�4�6<�e����g��nӿ���/\�rh�C���W��^r�����6��@e� ���B�D6c�z�0��(
Y�
���� pݬf/����Ry�a9�tr5c��>CJ���`o�6�ȐU?v�IL�Y��D�-A�&=WD� M��Q�pU)r�{�{

!��#�;���[7dN���mX��S�A�H��r���}Aľh!����
�;K�4���~2��	9��N7Q�vD>t����g�ea>�!�Έ��E'~"�x�>h��,u�h(1*ڂ3#�x^�r6�u�0�'�U��{�4�)"�Qߝ�tk��H��W_����� ֓�5�U��g��K�+�_4c���_�Ah�(1�V'��]UG��}����&!�gS��N<���@/��І���R���b��S��aJ��"�h�M�[`�6�s�*�{V$Je����tH�Җ	dC2dT��cnj�2���8�H��os���x�$�9GN��Kl��𢡊B���C��R �x��0׃�4F��u�)���mH�~��e��m��|�y��	�*��>YFF+�6>H��-��N�/����~+$ǵ��x��f��Py�ڏi�5ȄBTr�t�.�p@1� l�NY����\�9�'�h��m�22^�u�y�U�^��*D<.�6�\�Q���c�i�<��&x�Ω��gMT��\�p�V# ��;L_AQ��؎�4�C�5j�K}���U����=;�A��H��+���T����v���>�gBm+J����^�d�ᎇ�������.·���`�}��#��m�M(��92�"\,;K逎�!��̙�'�k�I�׻5Fn��bTݲ��D��"�iz���z�L�-�9�rfF����~�
�S�<b����=��Z��<�4�T����[�-���DT�3B(����K��.m����|�\
j����0�\`��t�������C�Aa��>�+�6/��,4^�����*��� ���}��}d;&�����xJ�ء.-�sx�.B��N(�~#U�>���}�a}���x�7g"Bh���+S&��P�Χa�{�\�w#۬A����Xc[����X445'O���>:��j�4h�A�D]J�E�	=%ƅ��t�{D��]m`W<_��K|��-�<�I�u*��.1�C��)x�Ia���Ȝ��Bn^�6`�je�x�N��r;���\����"�	�1��_�⓵�kZ4?!".S��
L��h3D�⓬TcbD)��N�YY�"Q<�D��AwM��A2j���J7eKbX$"ǋ��Ί�>�D��V�v���(=���d�P���o�նP^��ߘ��zd\�⏅���n���^�6����緺if�Y��,�/5M$̭|S�.�V�<�H^ؐKd��c�hր��c��((s� \��S�EWƌGi��7H����FP���]�Z��Hc,J!c���WD�y�nm�X���o*E��6LH� ����]u�qˑN�5=�i��'����Z��w	φ|��
oK8�v�$�[��7�_��C��2�;Q[u�
i�	8<����b���ⲝ���Q��v�n9�6�K(��\>���(���Ǭ������;h�ӡT��00�[<�t.�C�P�s�l�ǀ�(��.;��.�.ׂ�f��P��F�_K,a�W���Z����gx;����3�O-!Rl�ݑ��@X�k��L7���Sj��:^"W<�.��A_oŬM���u�S_���I�E{�vI�IyI�����3�I�C��.�-H��R'��/��誧>猎�J�f�ڌ��X�|�)ڛjb&�"�zJǼ�Tm��8"�$6{��E�g$�a___7h1(� Em~�6Qlh�-\v��ǌ��� �ֹ�!n@0��D����B��Rï�0�Z� 34�+J4q�.��s���GjJ���7��6�`}�Ay�>���	;�����^�ʶ��%��bE��&��p�|����J����r�|�܁�*^)We6�!� W��i�S���������/ ��9���I��:���:E� cu=�}�2�;E7��2��/8��PTB_���r)@[����y/����H�vA�6�u��8GnБ�$�5,=m��� ��P�M|��܋�a>��ȗ�d��`!�
���i+�C����z���!���>������R���Ĉ�e	��e,���Q��@\\\Q
�N, .LI���r5ǒ�?h�N����/?�6�5�������glb��p� pp`��;� ��~Ӓ)��/k՜�I���\4J1+��t�>���->C�6�x��qq�3qy�ձ,�GP�Ğ�/?}F䳔O����赎Od��>P>��p�d�E�-i"��t��W��D��7q3sWL��4�
J����S���H0�Y�����RL�FzĻz��P�9�-Xh��sҷ2�L�a}��r$��(����o@�t$:}vVe��v3��̚$����6wn�Z#�Us�����S��bz9�b��rԉ]H�`^C�������n�I\� ez��
����Es���E��3�Ǐ����I��nb�1(��'�W�:4�Q���2��5��5(W5����}���K�	�gn�"ӡ���gj�f
�rW;���ئXˎ+)����@]{�>I�=a=oh��sà��~���D���k�Q��et�&��'M�����ܷHj��߼Ÿ�7�z
�qLIŜV�8��d��f�F����!/�'�v�x�0�9V:�n�0�(y���(R��N_z��i�:7qziV�Eņ;E�D���F�SP���)g���(y�O��ys���;Ґ�= 3��V�a�����26is�J�11ty�٪�NvNl�S��w�	eV����J4x[[������Q�kj[D���}B��T�^v���Z����f�_i{%:�dj�(���,T��D*c�n�{�Vs ��߀s�q& �ɻS:�*��B��iuy_�!3r���Շ��_�^rqZV$+Ж\����7un��M ��@�����E��G��VhE[��-�q\VQ�=[EE���I���������4�d�i�|
ǯ E�sp"M*LzXn6��l߄l�_4��Li��.0�'��_,;�<��7z�ƚ�{�"�f}rFg��F'�/~��" }w��>-%�Y�慽u�9�A����6<�� k~o$/c�:t�@Y��zеԏ5ۉ˪���R]�ۍ�����[�l<I\t{٨V��{3.n��"8���"�d�Q���������$�4��)����%�)��i��z���Y���ϯb�4���+��I���k�JWĺ/p
�X��m��>���3s�XdY��s�"���xן������/��ײ�b律ⴵ&� ��ZB[��_7[��ˉ�'���Q??��������d/(�u�,{{���R�(BHӽaB^GN.�T�������-X�P����Ai���0��6�D�ӭG�dH~�Lfʇ%J��䛬D����`��`�KVQ�w��;��|y�������L�u��1�9��P��P������䀹i[���-s��S����I��������y���C��e.K�tkϓ#"��.�՜O�x���I����]��KPbӜ���#GrCo��.��@�H�~\cZ�� *)Ɩ,��-����^���:sI؟q�UQ��d
�V/�����c�M�V�tc������jv�}��r_�c��Vp��ag�-C�&%?낌�2ΞQחQ4|BD?F�s��ζY.���K?�x��~�$	�MZ�I˧?�I�Fm��y�����Ͷ-�z����\l/�ԁj�J���7�jS�7��_C�F��4�d��֒!��ۜ]?�������|J�5w��A��Ľ���nH 4��/3������ ���	h?/�X?��q�y[�g1�s���+�b���\��R]� �p�_3S4�����|�`��6Y�/�Vp�K��~d+�]O����'�|�VW�d����=×�DU����>G
Y��d�tYsb�I	�OO�V�I4B1�QJ�"߂����}�)����� ��b!����1�/v��"4�3T����dn�7`��"T��kj��ͧ�6dY�V�N�鿇(h�Z���a��P�#���N{��&�X��lL̝�izw��^���g�т5I]���r)P���j�EJ�{8q���O��{���i�Ґ��Ldg�L�!��z9���3I�S�͡�!�Lm���+�V��C��/�zsǩ��H�n���xr��W�44�Ox!���c���P�4�7w�N0�	բ����l#�?��+�[�]������r�:HVXۮ'q��j��#�:���F�����Q�ݽ��g.���8�~)i�Mԅ���{.Od�	�F��ͮ/�� $�
��Z����Cd����I��v�՘�d�P.Rq�n`�����9y���-b!���L�Q2�𬍫7��z�&XL�lҢ���͛-j-s��TfNaaaZ��?]���\�;��VZ����=\��b@d��[���[��O{6p&�3|DJ�$��'C���o��c�8��E\�*-j�}ٶ^�7�)Z�k:�]��G�"{�bּR�6]�w�%�e�F@�~��ږ#�k={e^{��M佃�]�O��b��ݍ���G���xKP����]e�n?�D�v�J-�G*��H޿���C�'��	��F�&kE�wT���5�Q��ӱ�]�Hjz6�<6�ҁHT[/0;�5'����')�i3�ޛDQ��0���i ���"�p��\R�ս1��=a,#�eVw���+�ߑE�U7)�6�Ns.�1M���y��&g�ScHݟxm^�v"�囧c����1�W_�;q���I7�秤 �e�0�. ��!��̀,Ϩo/()�<��o�@$u5��e�=�L��[������3��"������5��hTD���T���[�#���b��R.�6�}����܇C�d*���y2�S�f�b}��F^��g&�_Ify�\���Ə��b�a/(��͏�m�3X�qN��h��w�9?�z+r��$�T�l�&y��ȘP�`ˎ�#�7�Uo�����^��Z= �3�%�ۥ��ѣ�T�H�;��~�M0���?gL���#I5mK�
�h}�c��+�ε�w/������kg��'��h@����h�VE��jW�B���X*9���6̹�^�E^]�GMH5�k���r�<Sg�BRS����\>V5� =������͊���͙
�%�S��������y��EÚ�����4<îs^�sB�;�O]b�i��#����tΌ$կn�����Z��8�39C��\1QrV�F�&���(�D5�	F�̇�{<�I@luK{��RpD���d�C(m��1@��jD5�zq!��q�
wD�~,]U�+���w~Ո�R{�9jο3�3F^�G��_��S	�׌<�T��_*�9W1ƍK�t�l#.���3�%S���]���äΥϳtJ��+�ڟ�fA�9��.��ƶ=�X��a[��b�0��.��1icZv�=4'U��,�&MΪ�\5�����T$iX��齦�II^~�:��	��?�4����������n�܎�JY狐���E������ ��'�_m�)ɓ_�@�&��!��A�w����Zh�m�TzB)\J'EL�*-k"'��ɽ�������kH���(���j���<�'mZ0\oh���?��lI4�����s��&p�O�K�鄅|aW_~�:$�B��=Yfz��c�W{�z&(�݃\妡���c��v�֘��HA�M�E���݊JI��ʧp��f �C��j�z��GoN0��$y���2e_���w�r_(�:�`M���^~��q��u|u�����.���2�;d�v8���D: ��\| pV�x�=qm���'[[�LC��E�Y�ԓ�����9WI�������|�������1��Qf�}�s�1�M��W�B~��n����y��>O�W��{c�h��f"���"=�$U�J��76=`�ѱ�^^<���7���K�jo��p��N���@j_%��R/a����ݤ:�w��=y�ş��;�-��h�F�0��� ^^=i�W� <��_OZlE����Ɠz�o�ym����ɚ�X�o�o�U�u:�E��*�j����2���[v������h&Y�br;}�K��a�?�.�F��F�<)��ꆚOUj�
�T��F`�G��b�X�'RIqX���䥟w���z������|�ΗG��� Vhc8-vo)Y��R�P�C� �Ԏ�����������Tְ�Z�ɢ��e=!,S|��g��|5%��t��c�fr��(������9�?�*���dpKs�4��_R��F>��z|2�2Պ��ɾV���G�����!��m�:����0�C�򷏯���[��,-�W{��垭IQ��ꬨRM�D�wW��6�i����mq_�o[����\30`rt���.��"G��$��w6xl��&�������?a.�,Rk0���Z���)�r|�ț�H�"���5��C��̀��/?���l�GY�al�u?t�=4s��W���7����?B\��'%�D䔶�,$�Ψ��ۘ%��0�"�f�C�P<��~VG��F7������*��oE@��>M��q��R��mR���E\~�Q\ET���q�����`C���RSW���>S ͹#����<59z��#^�e���ڒ���2�SXJK"�6�9L��|=����hH��3�k��%���\^m�>Q��RF�&ҕդ���~?	!���k�?�H�(���/��x¿�mˋ;������ |o�U**���?>���A����nw�s\a���������f ��u�Tqc�����	0�U��Py��6F���Z���ړ�"��R�%�Q����׃���))� >��:��_����A2����n��u��E��|6�����f�.y�����E�ʿ�-�$=V\cmRJA:�U>x:�bɘ�\��UZ�T
ō��;� ޤ%ݸ�<���i*BR�bJ��-�'q���l]d*��;�5C[�D����$�C�ҁ+�o���&�0�1�M򿙙�b�!��8ȝ�_Sd5���^X���)���8���^K�k6����Yb�;7tU3o���Q��1�G����b�i�@��.Ss�`��*���f�B(����>�mX�8M��-r�����,�c6�}���*��MXwJ����9x��7�� � ��7j"�Ú���st��P*n9�B&6�)s8� ��ǧ��
�\]T�%�16f����S�7=����lT�L��h���m�y��ƩfΔ#��U�%�lip�)�S'���o��9��y�����)�z���0-ȥ�W)��[�ѷ2���9ØB!{��t*�HϺ$M��zu�Cv6��=֨����{��J�`c��f�,�'�u|o��6dFv;�y>�5 8�O�-���6=���؋������=�6Rn[#�R��ߥ��t���Ly���7v����=3�9�g��,]�@u4�d�t
��4�g?��K��
Ƚ����?|�P{�
DnD�� U*���0������!ޑX�֪�-�"�v�o�Sy{��B�p�fE��_��K*)����� hej�l���}t���:��j�]����C7��w ���@ͥ��Y fRf��3Mv�K�;[�M	c��6&O��4zaa-�%-��Ĕ^�B�?��N��<cH3�,���'ͼ �������u�b��pE\�����ƺ�����,���|�v�IGn"-xV+h�&�s�.�&Ś,t�B�������L��v@m���o���'��U�oN����~�*�����$}��@�:��7"#�v�����q4q��0.L!�ܖ���tNZ���YI|�̣�PԒ6�����w�}��ݚy�yC1�w/� mP�ܓ�;)��ܙ���t�ӫ���� <+�@�bm<��^sZ8{l('�,��sڧ�p����1a���Q)�踁�-*��K-��,��R��2��b�,h¬��`rAH	��[�ҙ���3�-8���	@߫
!�Q�uv�T����j����B�-�$l5�]GN�$����A���&=s���VD���)wܥ�8���q�;��X
��E����ωEĥ���@Mo!��m9I��1Y��$t�b�o�����E�M�al;P��C";���� U�C�:��|��pa�HB���0��FM=�l ����jF�u�uZ�,��vi���p�9��0�����%z�����4�3��`O��P��g��zL����Qt&�ET�Ĭ2TN*d�I��Y?��	�b!��ͭCW(�K�0��Z-�����~� ֲdyV�:����V(�|�%�~��V8��If�y����������S,�����`�����?M��~0��d$���a� ��4-�9y&���=4a�}N �(d������Nv�^����b�C���񎬟����������	�\���vkŜ������H�Ǆ�=�����~�9�Sh;�V��J����&j?_a��8�Ø�% E��(��`YP��B}L^�NEg&�nc�V��Q\m�R�ŷT���	���E�?����L�(�>L{���R��΄������+m�6���d��ɦ�<dz����Fؐk��
�^��������s�:�Ҟ�+0���z��d-��n�n�Ie��*e�
�K���u$m����.� �q���^7&�����#Y��I\��Z!L��u�5cL�/��]̝��<� ��wi�H}e
e��n��_��+�%!)��[� ��dٍ�SF��Gɿ�9o.�>��c$|٭!/S��]�F��*vC�JI�	�صk�VQS��*����HܸS�p�|oBߨN�P�M.����p�fj����Z����3DP��0����ʓ�w�U��#��V�����B�%�G��+*���,
οπ�O���G%�A^j�׋vb6�H�/9���k}��jna�њ)�9��./#c�5��&M\Lt���96g�QaJ
L��%�^��!8�龘ZB�g���GB�%�9�{��κ�Hբ���8ti��%A�|9=�<��>s�6�ן� 6M�ⴲD���s`�YQ�����c�^��dOk��v�i���&_�OnZ�.SrbᦹFލ�$']��Al�@!���ǡ���봜������FV�'��������0/�w��"o����ڼyϳW|M��5s8m[��ɾPen諔�(&�K;i4L4��L�,������J~���M6��i�֧����}�Y�3�dV1 o���u����]!q�� �j.Tg=���=��d��p���g���1w���?NhU�l�����ќ�L�H����ڌ4�kϡˁ&��7�B�s8�@O��ّFޯ��:� =�-���:�z�$ɼ\��d��D_���B�Ml��%�r�'{�ԣfL�
�Y���K��NHRc#�2�ˡ���0����xtm朖����H�l~�|���p���IQ�r"S���N"�A~���i���oa�8�qz���p�͌���]fZ��1��.���d��gn���)d��Xa\ߤe��&a�L��"A�փFB �[�sda{�k����uЈ q`eG��VM���FQ�Fu��C�b��Έ�VFZή�bw_����e��M�"��e�;PZ�E��j�}��+�'W�-�J��
b1�[5#oK=�,#��*������+1�jzV�G����}��O��,+�%3���fŞu�����1ov���x�x�8p�������nV>��Q7#��89����]cX?eSw}��F�/��l�er']N�\�m������r�	B�7�F��q:EW��͛�]o���06�*Rb��,��iz��=_ZG�G�ٕ���N�޹�Ĝ�I�^�5�(l�a, rK�ø.����о�FZt��j��;%��p���]�ts�27nt�,����
V����:�m��*����F�@,]7����}u�����j;�]���m׆��Ɉrl�QU�����O����o]T
6�j�49Wd6;�Q�J�?�.{�Ű�+�Sjˠ �/�/��?&j,&��W����6i�E���s�X�ŀ�9sg<����S�Ӂ�����F���/���Qc��v��R���}�����g#�8tk�$����f��8"�r@�>'<��;�u�@pC�@�^�
�K�ls�(����$������M�,T��ϰ�zϲ�ȇ��L���ƀ;b���%�g��Y���f�]��[Q�-��1�U�EQL6��(�թfU���T���\kdb��ͻ���LS(J)5�w���J���n����6M!�=��w�#Y����j����^��?�:J�a7���e0�m�H����{�R�����f��;S*���ef�����?��	���75 s�x_c�ݯ���>�G�;Oy#��|F��j�lf�{�ύ���puˉd\�lSwǋ��I�����"RF�/6�F��ps|��d��#i��H��-���DGq�����Q�JN%�L;�S����ڔ�%ǣ�+,6��:���w	��E������?R`����%�c�uĀ��+N6�4��9�T�������7�V�_5Vo>,"���2�ߘ�N�������"�SQ\��N�MV�LrG��/�Ͳ"WS䂀+���by/�T��=;��Ks��m����t�-6z���7?�e$�����/���>E_�k������5���}j@�������A߉E=�X'����j2442�I��I##����a#�<-<M���l��F���'g&�F Q������O.Pi�^�)Mut�A��޾L(_�kV���ylyF�qi���<=-�O�R�/�U)&F�����$u��x��Ɣ,����0��R�v#��CϘ���`�xJщ.��RO_��N��V 0���2��dY��Vj�ڥ��������+��j���R�ȭPYn�'d*S�.�[�R�&���=���P��ص�cOc��dP_Y����e,��93����?^�s���|>�����<�9g2_W�2CB�l8�o �]��b|�9�zŠZ;�'�hͻj/���3�~��^[ ��N��.B���Y6b��̥|�8�S���&ùd
U\�%��bE�D*�c���M?֏ B�X��)-�0���M�Ȭ��;�ڙT�J�d"7����jޯ��S]�w1�GG:���)?�2]�*��������`I@�лf���+[�<��B)���ܢ����Q�r^+j"�𷠹Xm���(��$!�+bI)������(j�k���46w�_�B��A��r�\d�q��Q?&�s �6��n��D4��Q�Ws)1��X'򤨅�+�
8t�[ӫ�SXb���������@UX'5�w0C�p�G А�ZE*F�������a]� ������^��q��p�.���	����6o��D[B�m�掉Y���k���5�z0uM���9eG��H�a��l���ޥ��j����a���'do�R?_���˾T ��韜{�OV���TM%C�(���x�ݰ6�$Ѓ�Z{��8�(�>�ܨ�Li��jP��[}�r�Pڸ���;/�,]��>Fn��
��?����_"��
H�f��?_�~*Ew�fFa�1����L�U�8���I�R=R�1@k������S�׹�?J
Lj-G�������������Z�:���FB�0� ������2TZ�փ�i���s��.KͿ.%fS��\~ig�\� �[���n�Yx��$�3��m�& ��D&C\M����f��|�)wZ;�a�Y\:/����ї��f�x�X�+�i����B����N�z��1{ �_���w�8��0�ެ�#�A�L��g����.�տ4j�oٔ1�u>��|���ɧ�e�?�kdeK	i��֪Ň���0%礴V��P��Ai�:rQ�?��hX-YC~�
Z4b�����2�)	o+(i��|��a�e0�<]��c}U�8o��\c>Wؼ ��oh�t �|�	���O)Fc3瀫�}+���,C�V���]�6pV�Tc�E2o���a�֭Y�$�t���/�l����'�ᗀ�S��ѶoX5Av�����ǒ᪷���?�\�� �F�j5���3r�!����"�#V<�\c�����X�\�gN]�V� ���s�����tpV��Ӫ�%�\շ��[N���(t쿙A,A�y�h>,֣��*4��1
�?����!$-3����xP�~a~�&΢��#����pb��q��3�N��f�����9}��<��DKA��(��]\j�����!��ak�]BL^�z ����CQ9SCg^���<�7�J�H�=��|4��,��d��� ��7�գ�Μ�y�u�J?1�`L�M��=&_F�2����\TV���Z�\Yˀ��A��j�9��9e�"8[�Y �D�M���f��`�:}Z��Wr|lq�$)���s2�φ@�n,���R�$N,sѓ�@�4e�E�??����*
|r*G_mīڇ���꒙�t��	���M���<�ɪ�f�jf��&��Cq�z,#M�0cMd0��P�%�4i���O�	�A+á���@����O�0�@����gA�}�������Z��s�a�$k�'��vJ~c���rݵ����DK�|�]v����d�� ��@���9[�"�0��S�|=�. ˑZ�pM��(szq�.�F:�\�&2��EZR�-�,���$�?H�SǀS�"�M�\��6��!�)�E��5a�L0���u��t�įP6F�
=bw�� �m0�~�-���ڧZ8���v0��w������@i��~z��se���J=Ȇ������, T_җd���Ϝ�MцCndH��#�Cm�V��)�>��dU`x&��{G���g/��E3�f3�D�$�9xڬ���F�Zm貦.O���	�b}
3�km@`��DG[�$x���#$����y�P�E�[8��Z�_�|��b���-
��`}1ZC���aH<������F3�Y�_W^<��rȚ�JK���m?��6�_%_��6��Q,w`o��l���6b�x�:�y(�G�2�q�U�l��u$����|�:Փ�Ű �(��U��$NS��+���]��N�XNX�k��9�d�a�=}���tvB%6C߰�B��0`�9lr��#-��[�b����x�(#g����=�m����k����s�/!��9 p��t'��d�7-�2�6j�!���
�#{5��ĕe����O�G?��4Aƥ޶pF�߲r�3�9�E_���@A��0c�-����(��=����oQ�ɩwJ�{+y'yAAJ�Z�Yz�~��K@�@���{fЄ=&g���3�~��Ф�\5��uk���h�G©>Y'�Ճ�=?&��)�D���.�(-�{�Y�? �2�`����k�3�q��Dӟ��|vs�gx�)|l�� } ��������-]7��,G��G܇�MY ;r�l��כhEb|;�b�\����)!��jKoZ��O?�u(9`�o���w�J{��_���La���CO�r�g���뫺9m�� ���K ���|d�ˈȴ���}����4�ǋ�vEU�FNj�U}S$9�(����Yf��v�_$Y�&����2c�׭?�/ k���:�{�K�k��S	�H��=	�8�w���B  �h����b���'M�*YK}U�B)����z̆�	4@�#Q�M \}�r�غ�]�W��!-�ӥ?9i�	\Gn���s%�X�M�}RV���6#	�)��0�X��Db�M�eΠ�*��� ��xr�����ksx�id�����K�j��;���Aw�i�=��9����^�7+��ٖț��Ҷ#����P�3��B��?_~��4X�;��k�H��D@�q �� �:�UVN �a�M�23�6IS35����ֆ���W��%���\���
�V�Y� �Z��YN���Y�!�l��쫵��D���[@�-V!��H)�J��YZ۷V-��ؐ3l��̩���V�,4�P������0�C>�Ӿ	��$`#wP=�cy���
�-��۰���澯wҦ�?9�S$����p���%jb�У�K�Z�͋����G�{�r�g#X�d!�7��$0�D���KK��]����7�,�� ��<��O]�>�p�`��.9q~e�L�+)��B��O��z�����>${�ݪ��rĦ�}�:�iZ��X5"fK��2�n�oWz^h�Ð�t�
v+��	��9C�{��Z	��	6�/����7:϶d�BGc1'�p.݄Ο�n�]�[���*?A�dx�����8�LT�@<��i����f��H_������$rIx�1��k��Vh��#�<�@��{�8��}�����(S�qp?�(ѕÒJb��}sף�F�8&��E`B>
�i�^1�K���a����S�?8���t�u2�M��"�z@�_�� j7,n�t����$�t)Rq��9";�2��[;Y#����i``��^�<g�R�2K��	�<�y
K�G�E��u��~� ��i��61u��:�v���ם�r�D��[��/l� ����b���+�'���d�n���}H��1)FTׁ��<�FQ?{��i�����g0����� y��f���pW��<�P_C,(_7�·�SY����\���	�{q�}X�
����!�kabͺ���v s�Ь. \�ՙn+�kJ����
���;1��X�vԎ��\�M�4�`?�El�wW-(:��T�?A"�m�������6�ΐ��.�{�y^��d�$m)<���bV�n�����W�t������#R�
zu����,��,���1ޕu0��l[@d4=�h����z���P�i��e)���;G��at��^[m��cW�kq��mZ^蝄�<b��t����\4�G�y�Z��b������*uy[�Y��?K�DS"���P�eM��>.��oV�Ꙁ+�H��i*��@��ϔ=��B�q��<��I�v֗��:g-��y*���U[k>�.�V��̑�]��U{X�> ϱw�.~��ŗ�2����E�.N��Jv\���(��5mn�T?	��b`�&D P����Ta�Ȕ��^��Z8DՂ����^��ΡT����:3LxG��g���Y�~SB�P
��p1��w�sL���i��5�> ����J��/QM}������Mln�-������o��b��D���������Җۄ���J1�91�&/�S
�Y�·[;���j+����C���t�cz� S���.�����Q�%|�z�@WV��~C�œ��!NC��0�GY!�C^��_K�a�]�� ��*��J�3�R)>=�,>�s��a��6��f��ne��0G��(�^� Xc3��Hb=��Nd?��+��"�Z��Sr2���ć�q,xB�!���38�.�R-I�-(���g��4_*R���S�����Ю[��=K$p���eBa�)7�\(n���o�i���hi^�ILN�)@>��z��~k�2�����U/B�4�@.�'��˖8��$]���� �PIt���V�9���~������NΊ�LU��I[*�SN�K��N�C �j��N h#f�FL�Edi9���ޥ
˨:�@��ҭ�j�fj�S���B.����6��ץul������b��76x��r��P~.zL���A+ٛ���/e�_�U�綱p����\9V�Ҝ���4�m'\�%u����'���!o/j\����ÿoy���^My��G_d8h;�o���-���"ʚ8����'�&T�&�MI��9��`�ޡ�%ʸт�S��>��bE��;�C>����1�d2V�=.|4�-f�\� &�xʕ$��D�N|�����*�zj��?l`�~�Z��EȜi�/�� '^�;H��Eќ��/�UZ���7S�S�����{�ظh���Q�����˫1��}���K\��?�,�:*eM��!-R�%�nW2[�!���������B��T�yl� -��e�-��m��瑚Ѷ�UCh�
�3&�Cv~W�E_���ު񱓸��cp��.É�� �b��r�}�,�V�7�~WYխNei�]��ӣ:�lI&�X�J������ǵmЇ��;A��<�.��Q����Yd�:�
�%3��m@�yCغ7��㧱��2��lCC���R`V�w����BB�9�􀇗χ�`���՞�g=��kxn}᪤|t�Y����dAvI���g�ݮ�*h��
�7�>X$�3ະ8P��vi��(�LK�����ھ���W\F8��p�Np#��AwC��sĴ��j����q�I�E��:z�>����FHb�n�GS��y�E�R�t�J����O���Zb����p�Y ��o�7՟���yr�p 8�)�p�$��3���N�a�~z?����K�-��������x�w��V������񌚼�.����f����PK�X* ��0jwA��b��
M�C�J������3ป�*.�Y0oY@�u�٠�4��$X���G'��Y{(⋢:p��3%�^��Nf�v�z�P��A��"�l'lE�;��Jē��|s)��\��9n���_f^$zs�G,߽d�hR�9$�3��Ch���-���-�����gb�a�K�eee���d��ץd`��[�I;��`� �}O� ��HFx{f��\�\-'���k�佷�x��0^�#�ֆB�vtt\���v�x�4�W���F\���j���k"HST�	���\M$���~��vq�+%w?[a��d��%V9w(m;B��/�Q9D���YfU$yi�eX���hP$è����ג⊊�fX$��V:Û򂮜����<P�
�,G�/`q	|�̟��~X�,�JL��rA��چ������J|b
m��H�e���t ��K���?��6��~�K���3�@+)��f��%��G�C{�A���$sd�]f�%]JJ�R�SOi��q�ȇq�!��qP�i�_���ȼ��h���88���-28��z�6b���+�XB �ўJ��͒>�w1��e����q� 7�wZ�e��)P+STTb�����Ҕ� ��.쬝΢0�߈qUڝ�2r ���Ӏ�]��@	�l��\��~�,��k�M�;7db�kZZZػҟ�.Nld+�3r �Y�_�R��>� ��ޗҳ>i���V��Va�1D�E0�kϭ��a�����EC� 4���DE�A#奂v�J�a�ڤ�U�3����x�К"���rに�srk͈����y�P�aH}k3π��S��
���{E'��t��_C�Q�g]9�\J`��G�ť��lL����r%,�9U�����͏����U�M�]��#�1܆ϓ�8���6�:�FM���@�Ȧ��K���>��7,��?Ö�,�1��[OU+VN�)?�$p.�q,��U������P�����,�9�������:��E)�N[��=�K�|��C��uL#,�����z�f� ]�PФI�0�']�ʹ�e�g��z=;�ٸ��Z QhB/i���<{����������hd��0����9�����*辪�j�ӏ�|1���Ɗ��T��� �k�Mi�z9]K��}πG�RR7�	�㭹����ˮC3��άUY�%� ��)���;ef]b�?���2	�����6A�����>*%+�֍�j|�y��Hܣ>)�3�Pf%��JSo�~T� <�=W���j,`�Q��� "E��(˅8�`bb��3޶w��J�6���c`��^?^�);qV`]�;���M�p"�� ��[��@���ʡ!{~�;	�:�/l�{䇟�[�Z���Es=_���{�=�րᯏ�zP?�SA��d�*�>��"[�7�^��%=�<D���k�������"� �[��%�Ƭb[�,�7��U~s
�P2K9[}V�wƛ���+�6�M���+2�|��M�ڵoƊ��4K����IY��X�P�|���Cc|m\��2��5Rzn<1�/:_�(A�AN����K5�r���z�#e��b���\Ȉ�]�fK����a)ω�iLi�Iݦ�Ȩ����Y����n��4?��U�5d���N�W��UĞ��&'�p�+��D�GC� ��q
i�%F���ٰ�z6�'���B5�Ĺ5��W�3԰�,h�w��e�c~'�����"_1��.�'�����	�
�^к��c��d����OQ)Y��sb"��7�Ŏ7���Sn� $���e�yVh���IÔL�����(8l,w��X�ΗF��u
���q@NG�w!�g����l�z��^O�3�{c�<�N}�e!�U"�nZ� �giK��1Il:o��3K���Ok�=C�آ~¼ҾT�8f�:�M�(z�mL�� ��bJ$�$u�`��M���Q�g�k���2�g[��6�ǥ�2��p��[���%&����w~�B{=�&-��N��f���Y�m��s��$a������x]����(z	_���jϙ�:����BM��-n�I��#�G�`�6�z ��f��؜������(��.��1 ���Ng䅣�3G�D��A���'1��Ǔ�'���
iU�YJO@Z�נ�*��,�X.�MR����=6�f/o]P���8K,;�����H���=87ϓ�48��d3�
�\Z��V�E��<���Ѡ.����5SWF�՛�ڋ���oa6ܨ������ނ�ٮ�M���?E��Oʭ��0{o��:A(�O�*[���7_��,X��DȧB�w`H�K�R7ΰ�����m�f�ΐFjir_h��w��.�����=���TjZ���%�)�)١�����kJ]|=v$�"�t�.�B���(�d6�q�ɦ�0�'_��[�X�����k	��S1��n}W�X�֐���>��ڑ�W6��K!H�x�N��|��̰�jf����q�C�`����w8vSQ1]��+J4����:�^� @B��xX�>�O��8,B
89�nS;i���k8V~���[P�GGG�0��Č��a�E�<b=h�$���>E1$�%[��s�S�v���}q�5��܈�J�R�ܐ���$��e"H�-Ѵ�5�!�~����*}~��F��(9RӔ%���!��.�VT)`��_�V�����/I�7�b��a@�;o�?V���<���������l�Ѥm�1&�~`idd$�*iP&�E�cAJ�����U�<����� �`��tZ���z�U�8�Ջ^����/�=�	<˩x��T3 ��N�k���G�^�_kB{z�h�FD ����~��,���A[̈́s��J죀YX�pa�Z���U���d�N-l½a݆���7$�B��'v$����x�!��Hn�If>���Xgs��%o}��"p� �,2=5��s���s�%�)�#�rW��Q�����z��)�b�Y��>x>Z)��7G�y{F�ft��złA���BP2bޒY���& ����@���$Y��r�	���V|��F�n%��B��t��$@#��#-���0���v�?=��c*q7S��=��qR���O ��n�X��ϮZ
 8/���j�k�`��!���Ub�:�ښ��TOϜ��+���SF�.���.�a��(H���+�~�9M�7�Y�BMRRU3�Dce�>�RRcaշ/��봣����N�r4,���D���><�l#��9�Ÿ�]�4���T˘����
y{��T��>���/Q]���F�-B.B�NSKl�DP��`C� �ч@l��ǳGǹ��}��齾3zL����{��>E�}q�,53��y"���3\=���������x�A�}c��?�k{�s�ob�f����
'�#�%���b��7㑟�^>!��PS�j4|^d���Ic�J�@�x�L�����<�0���j�Q��5��^`H�MQ&��4�!����O���"�ow��4���q�e��m=�aV���W��$z��<�.&�UJ"iOVti�/�����8?�1�2�4�j�jW[��lDr�䀈`�1�/���&9%3IX�
簫�X��i�Y�qx��G����.�y`��g�{S�e�
Jr�5�>�#�җ�NƜ��2���'�
�(�u�;d�~����m�ˌ�b�	]}�!� ��t�ϗ9�9�gv28���Jf�r�����c�O���}u蠗t��!3^KH�os0?��*���Z���H�&=9tUFx��mUxj����j��j����kϮ¬����>�)@����Ƅ�s&+XL]�K��Ģ�\ϒ�F�ӏB
@�bN��Y�#e�pR��I'(��fr	ܛ�K��[yثT����d��}�lِ�O�x����3��;����888(�q���^�5��(*Z{�.Q��L��v�������F��@N؁f���\�%�|*v.���rD}�PɌfPH�{�Z�+��,��і�>���Ȱ�mmmOa�3�ᦑ����IGE,8�B�a��c&�ډՂ�:�\�H.�{F��%l�K\O�+���d��ؓ�Q�T�q���SlI����A�!ۤ�u,�"�˓Wr�;�a�^�,H��M�U(��ݰ��:�����F7>���&��ʿ@��L9
j;vBK����͢�cW�|��	���{�_�y��̜=pc��� �8���8o����%�`�f��{�����a܌�T�P�&�u?{����cb];�	�J,�X�����$��	��iry��.+*)�Sҽ�֠Rŉ���DX�7��pQ�J��$(a�-�r�>Q9�o�K��o�����BAk͵�� ���9��~Mj��R�D�S�4����ˬ����G��R��6)� ���5�����ƛ3����`<�V�u<3i,�ڵ�"خ�.�
��-��>W�ڤ�6ň&G�M	�g�M?�C~�U/I����Gy"웽۔i�;��wן�L���Tg+��A������UMu������f/�dH䣝��~�lE�9����d������I��ڧ�N�*�|�;[=c!J��x���	E'*PG��U�}���C%������k�%���j�)#e�SUS�x���y��Cu��'� . �0��;�fĥt���Z|����oR�mU��C��7"H��
X�exݞئ�J7��H����}G�᳣��a>�h��WD���i�@�����@�ދ�	x����kg2c�n���6�q���
z�������n���5?�wǙ�ҍX���W��V)��z�՘
,
���%�U��:���`fcס�l9a�j�5T`?
�W��+R�%�K �N��(]Wr�*W�]�Ӳ�<7�E�Ԝ������ �)�		eNa?�h����M6G��k}� ��n��pn�u��x:-o��ްc���B�d�Uw/�`�'�>#H��Wb�sJT穽sssE111j]���l���ۤղP�'}��������4`�,��{߬7���+m�<u�1��T��q���VH�?jP�̯�;z@�%E~f �V�+-��G���^�zT8��Drf�O��sF���'�D�Ϡ�߻<�}Ɨ&t5��x�I:Y�/�^綆>2�8�;4�i��ſ{����P͝l�\�(�˅�/%�� �
pA<�����p���&j�x��˫�!��&J�q���.o��.t,]Xdu�?�w�*h��Q�[�����3[�N���a��w�w�sm���ܴH�k���4fc����9��Їq��1�S׀㚺��|� s��\BdK<_I̟��F?��r8u?8@.��]]�3����
ٌf��<���ޘ
�k����,�߼�ؙ�}[�e�G��ӗ���B�h��!ޛ���eH���;~R�9�%#A��|[�&q,j�~yр���w�|J�� ��������2
��bJ�u��;���>��=?�{	�oW����
������^�o���G����08K4}M|���UPo �J�נ!cA��g׺Oչ�h��-��|���B�Qܓ�ځ���i������vx��m��I���*f|��D?1W~�W@5�vdr(jW1�E�=�k��s71�` ���D��D�|E��P��d����Q�$�j)�+ӗ�?ÚN>�:�,��H�<��v�w��.N,�H������Z��V�
yNOѽ�z��S�Ntc��x0@<H�J&%wYsEtf2��ۅ����dK�
)!^W�����	^�PF;�?�׳U=���m؏g��v�5�w�|A�����1d�*R_U����<�c8;�vCl�ގ�\�����o�H,M�`ŭH ��RF����:�N�!8reen����;sd/.���a�J�v%��� �w`,>�e�����y�Z�����@�G����N�H�2��Gy�(�
�!��Eu���e���3��0�.@SR���@������Fg��N*���$���}HO%|��W�NʜQc�� )����Ǐ�V�HZ�#�QO�1I��A�� M�M�O*�Y6��?VH��G�Jb� Z_�(J��'����n��G
[� 3/�j����;+	!�
[��B֟�:�%�}U��
�l3�f�*�(�|x�̋�Ê�y^A���'��P�?!�xy�(߁#}ԅ�2-D��c�X����$�>��r!��~ N�҇O�C@x�C�xͿ�g<ƀ�2K�x>�骽�(Yܹ�>��gb�^Y���0Ot6eWm�gس��u��잛\J��@M�1���
�M��д��*.�Uz�@�;Н��ff��pZw26�g�7���[��1�SR���j|B&������/��p"��*������//�g���x�K�+*sK�b{�y8NI)F����W�7��c�v��� н*�u�����r/`tw��;(2���hVkԩ|m��>�?��>E-��<�> �F�Qi�|�
v@�w���P6%2�B����;Mps���N�h���%Ǭ��r�ĆX<�#����\:�𽦀����='�ۄ��~0>E�Ja.�D�W���7��J8������G޲=@�wZjs���N_E�!bC^p��<�5J�L&S�{ei{@H�	�"�*��٫,�KX����h��Ő��̰_�M�Gu��>��1�)��NQ<PNޠ�c�"��y�xuwbt�UP3�ٔ\ӟ	�u C���0�ί[��i�����Rk���Z{�4������G��J��w�~:�f�����%.N$a����l���B$_�,�	XF��	Y�R`����(�� Wq���_�ʡ�K7!��N!����Sv�O�H�]�%,����`�&�xx�����F�B�(Ȅ4)���~��f�A˿Ïa��5ԷCP�S��2P�2`�Yj� ����G��j"�jR�|�ry)�\�"àEA*�,��
�} �����*S �*o�bO��� ��c����\[�߇!ͰS>�,�J�����W��Id�i��u^GH
^��?���$�m����4�՘�斸��N��k���!�5�m��'��81���Q?>4$��p�`��:��6�*!l}7�Qz��t����R����8��9�Y�P[�o�[Y9&I끯g�F�ID�_�SO w7͘������%�p\��!n�=>)���M�L��%�� >����C�����������Ѡ�������(��_��R@��3��r#;FC�gi�#
��P���o�}�j��"R%ol=�Qi��H!<&0ï������I..�h�CH )�֛��c�r��CJ=�luM.	��D�C�l�OL���,����Qw `P�.�ߧ�\v�5?��j?`����E�@�~���O~�ɲ�v4߽��֜eӆI�c��9,�A�7�G�������ܐ���S�Г8���OcE���ܹ��>� #������FA�� �QT���!g�D/h��Z�%�|6�9��6ZYA����K�����X5^���s�>���E׆�C�ۻ�A5�{�m�M:�W^R<:����8�����hE%dz&�%=��B���v2u3�i�TGa�9t"�;��4�L
��4V^�mA=d��п>�cA9t���N���2)��&�|L���y�.T��il[�����t�G1|�����5,]���s��x��b�!�sӻY�Dg��O�!d��E���!��o�烾vJ؆~��f���6ĝ:w�'�n���!����N��@^iL�&���UYޮ�E�/�*΢�ubo��n��Q���H�fd�t2!�8��������4L�.�V�xR����YEI�B.��8��C~3`�̾����R���RD��0�E�sֳ����y�Ri��Xj�mwOO����J�gC�@�؇��}�������i��_������f�׾~£�a����(����q3	� �z�1�l��J;x՞"{�o?1Qv�w�����	�+��8rs�n��+���5Un���M7!k���!<^���ċ��V�t1���,��YB9t�%>�D<|"OPG��s4Z(�PNC�PZ�;1��k��bib�߾�%�f2�����UI����Z[ZZ�:\� �:��4qK�V�-9RZ ��&,�;wN�|�����{�*�bBi�ӳ�=vt.��Sn�Jn_��F���M3N�1��
쏅=�T�����g�������v��u��Z�J�9%�p���	$�c���\������;|o����F���jY[[��?�^���fjb�pʫ*�{E���o��옷g����Y�'���O�.����}��0� �8�t����ɬ�X17��&��Q�,���R((�ɑ����O��eeKx$?4	�W���E;��{��pM��xm?�\����:��>�we܌�*�x��VVO��T0�	8y���\qbbbe.�o�> >��
��I'�;|�[�$�X0ϩ��k��z\JX(�ap�D���M�[��V��jqtҭ�oC��]K����������j��R��D%�4�À�sp`�א�7��\d�]SWw��j�%+�ؕ�q/Y0O	A�HP������OԷǥ���I�Hz�%��5�h���*~L�=�!�,�A��}�;~U���W�?m�
�����)�@��x_ �?=�-!E����'!6JY^A2�	���dX�R��!$��nD�O����a���}��0����ƃf�@Sj��x0Qk}5�QB��%j3kN1�R^\}�"�I�p`�� �*�@\��'���_��-)ᩘKo��$4` ; @&p���.�z��(��@���{���-�7�j���+:���ÇUٽpڜ�M�֜��`�N�-�j���d�Pj8� ��`�/��a̯�&�������fC"���J(w����������*y-����d�'�}y����@}��������7��ڡB���X��'*jI!80h���9�3�l���*��?@���K��*�q>~��0]�ꓭO�w	��΄7J�7<?���eO;����@��)Vu��m߫�[@����NS��U��;�4���%��.9%nO��)��&O2>����j�_�� ��]>�ܕ�M��T�q1����
�$�V �&�Ŝݞ����_<�;�;�)����jN+���M��7z���.N��V~P��哛Vs� %g�#J\���IpI�2�;�֎t��Z��-v;��}	>s��l�nHopXs�_�#�/�~)�����,or�'����m8鋟Y�i�����������y�ж��{�5��?�Nw�Q����-���h�v�p�_�Q��@�M��c��?��Pt+��\��������c�
�/i)ߍ���٥;�&������SJ/�MR�t	�7�WV����s��:��+pf���K��.�8_������|lg0�m����к�_-�7|�R�&�:�ۖ^+�TmSK=���H~��������\\�n+�Y���ĕ}LL;��S�t���]����L1���&V�hM`y�oʙQ�Wb�>˿�Nr��PcS�) ���]�)��s>�&.D���	�����i�.�Ja�4xݸ�Z�۷��o�O������ŷ��ʦܮG�>��0*�U�^g��a��n�:t�6(xk؁b�*�p��z��%��`�2��B���u-}��ZnzyW���O�5o����~��H*���N�s[��C��	
�ޝ�^�뵁���|��p��R������y��Z��o��w4&:z��䭖4�f�<hʣ�'�ݼW��[Fz�餯I����'�!=uHW��[I�c�g�mBI-����b&�/o�4����r�w%�q���w3����t�[`�⎬n��%�VH��N��J�{Y���O��6VD�(@z\���b�f��ү��o��K����@�F�����y8aSgI������R|��)�`�s��G���8�yr��y�9'��t�6���N�Mu^ʅ��;;�k�TYBm����vu���/V�oQ�D"�V��<�P2��4q����io���/-����þ�9���v��w��yn�̬�T�s4K�s���|]g��j��Э�;'�w�0�<Vz��)H7h���/��35��j�de�ZU�/�v8�o�w{$4b%/��i�;ׂyYd��+G:��y��碯��|#}�%�G`���w�v���<V2N���2����Mccc�U.�HV�W�k߱���{��T}�gaч��Q�kd쳯��K�-�����}�RK1�"����XA�D��q������N����|�tb��ܴW������9
�yTn�X���J�q��
k��@�?�pN����;l�h0�M�V��uv'�hQY�>�?�X��iz��%��?m}Bm���}"iT�����\��Y���2��Ƌ�'X������{1�Ҭ��fh��*�y��%�^XYYI}��G4���AX�랿�k;�Z�5޴ggx텈���r:�g�%�1-�e�r+��ǥ����h]xF*�]�4<�.+''�^�������ź�+�������L�W�K����+ߜ������>K�^+���h]���Ja �rr����<-sAeȁ�r���*m��XX�8���}n��%�F9`��c]�l����9�>�3���d2��VV��m� ����׾�nv���o^�M$�0��ٽ�r�L��Y����� �(�Fɱ9��	�륍�����5�=H%E��$ge�|�k��?�; doǏ�1����{�,��ݹs����>n���l5��󵶳��Sͪ����/�)?��>`y)�2~6�{��/�|V"_$��A�r׎)��P��am�yQ�7ͺjTq�䗄�A�w%���@��f��S��!=�N���B-�om�6n~&��Qf��k�w���;�Vs�� ��k����n���@���ҡ|R��o��{����_��]]������E�M�qi}���cx�]}�q[��� ���t��o��쾛���M �\��v�����`dd��������[䵛{}d�o�w���k��Φ�@��]�\c;�>�(TZu�]�j�O{���B�fE���M��7�#^��>�X�qǍNM9�z��������g�o��J�o,H�< w�색�j�b�B�%��P|Kw�gC���B�����	�RI�a�#�<_n���<���"��I�F���\\!�����5]�!�f�|nTh[���-96�Na��nUUT4�v��I�l���p���L%�l�����o�H�i�R�p;��oGt����F��v��wX �[z��'�_z�����)�G`��P?��i�X�x�j��v�f��U̥ٽ����uY�rRT@����V��\,]�t�]�qO�Y\Z(����n49��x�>/�7��y��0E�z�ݟ�?�-��0�~��]x����)@�q�Ϯ���vT8�]W����,�$�84���㲒�^y�h�6kI�ke�p�;o���#���a�4���k�Q�ht�����eSDˆ.����x��G��&�u��B7�P{��,&�[�B���0xpCCdܠ��B��w���#�ϥ�Hy4ix����Z�<옱��?�ˤj@A��GU�@��mHgxvtekG,�^Z�J����DO���׽��`�^F/�$^�T���A�۷�b�M��P5�ɰ���.������
�'�2~�Q<g�b���j�j��]��mz��|�KL7��0��Iކ�
oo<>7�X rɻ=I���{>��W��M���a����T�x��5����j��c0��ݝh $7z������_�-h~l���$];JU��q���6��"d�߁�;ݸ��}t���ڏ02�����O}Q��/���kl'%�;2�1��.F�w!���)��4�`���{aӞ����~�xg�.����`A��ۧ����:lJU��"����B-Л�k�p8�䉮=��ɋD��+r�x.���o���S�\��=���>G�Z��?���@�T�MP��;��]�m�?h�73H�~|����Ŷ�J���Ax�R����N;���7� ��_����r���c��zdjjb�<���a�X�Z�v���I)��{k��e�A#��3!&�
b�l���(���;R@@�`~����9�R �M���J�wנ�
�2�:���:?�N��%�S_�u��9|����U}�����>JL$v��4}��A��c��j�~}c��Yug�ȁ
0�~͵Ϧ�3��_�
cFGh��d�=<<*F�&����휦|�Q��e�[E��ϴ�Z.�*xʼw�����<�s�״�}V:^�D��s�I��'����`�"h-fp��{��c\��O4P���eL���D]�M�*��NM;����]>p����HOʣ~1��nĉ��W���]�J� �@��~�T��7�&P�?��E��͕)ߘ�y�V���A�c�r��#���U'�\CAѮ�^c������Ai��{����@����*@��_� �m��nRD�î�6IZWIX�yE��s�b�Z[U����@O��T�C`R.� � #�|�F�BDg��c���EGs��� ����������~P�&{{{#1�9�@�x�|wbk�m>iӞa��"ݠ)�r%���I�a���-X���4��;�Oϛ��͸�-�8a��3D����|���Lk��X��R։����\MMM?&��$eBr��$][���3bo����d�_-//�z�f�-��ǻ�{���e��K)���|�"\�H���\���5<��� )7n1>�ip��Ӷ�e�1
0��,�䭥����=���ǺUz����D4�v⻤ݜ�Z�	�B=��ȱ�1ء��i)=���(�0��UC�U��C�3���k�����56�"��*s:��+����m�`���EwF�����Ǘg�+W0t�h���E�=��C)����7�N�5>ǧREs��,;4~I��O�TI1y���tM�~����e���G�����%�T�m��P�H2�
�� T2mlIi24)2�d�2l��D���XGE		�mI�2��L�6Ŧ��?k��������w��:�w=�}�ϻ޵��^-BZR�A�LTD�mS;zyМ&,_�)L )�bHQD��I�;�Z�L�
��I�o�ԓ#��}��d�3�([8Jg|Qa~)���3��S��Ī�L&�vtx�b� ��t�D�/��́P|�G\��J�l:\9��>��߫��BJ򗩊_hƋ�����zf�<�P~�5x9��I&�`�#`W.x��,��8?��l�A����լ�p�;-j����u�6i�&n*��O�lL���m'o�)r�L�� �Mc���t�=�=[�t���M�'� �H�ڻ]�ˉ�������֕��$�h_����Ҩ��e�tF1,xc"�E#wH��B͵���i��3	�$�!w�+� ��
;5����o@�S���7㷼�͆G�w�%}y'��ۻr�@�^|��c�k�`���f>���餜����pP�Vvgs�
F������}�V��~�]�p��Z��X�2��/�e�uZT���q39��l�� #.	�'Źԟ>O��?�����hu��)�d��W��������z:\�nͲ�E�x�I$p�dWy��ŀ7�:���]���ng�B�o���=g��^�|Z������=�+7	Ġ���-���IH�����݌��ȓ���ӫ�e�
h5���I�ze�b�u�t����;�����ga��Y�H�����\�*�I�)��_�J�&}U�U=Z���IA���� ��q)"%��5�t��a5t�z���0�F$C��|8����Sy�-�o��*~�A� Ì���N�0t����E���~�Rė/C"�;�8�m�<�-5�vi��y�}��+U�K��3��a\�FkS>����~uA�`���˗��Xw�t��Uw��/���{Q�C�5\�k��Z�+g���&��O=������e1z!s���/������r��S��S��yk�l~ߌ���d��v�-�l��0���,;4��u�O�r{����h۳q
]Gw�����`F�V#/%�4_��!䜢���E&���dݦ�C;As�]$}wtt\�~��}�լ�:P�oϨ����U�y'���w��&�b ��.�1K	r|mQ��
������|�÷!����޾B$}�D�@k[��Н[̞�K�����*9��l��q�n�N�n�iL9�W��˅D���p���C�6�3�Y�OMg��t���5^�|7\\�AO��ݻW�-��jˉ5��_�.���f������u��,����w�x�*�̷fQ&J&K����J��	1�O��WO{s�pn�g����Iߔ5^��M���y:44������m|��c�u&'��Y:�A_����aV�x���i�����ȏ�#�*�m���wOVF��Fۖ����L���;���y;3�+,:�]�5���a����gO"����R��S�\�K��*^ tv"/7�\TL��J� Z�AR*����?n��D�teGU��ג�@�[�P*#�����5�Զ��ȓK��-yj�C�K�J(��	}�����B�����g&��q�NTWx_���pi[$3/���H�̩]WJ�u��?3��Z7��`�Q��3�EPy�x=s;����l���Ձ]J�Y/٩.���K��a�����]!�F
G}(��X���H��7��ţ�GM�VT�|s��ן?c��@�<#n�'������79��=�[I�LLLnCR�>-Ss.�����M�:p-YqH�Q`��v
�8�b�c�]�JMA�&�쒗��ҮO����p�V{G�b��-[����}��9|b~��#�r22���>p�U����H_�@����MW=�z��,�hZ�kr�+��n\��u�O�8��T*�MV��j?�� �+��)��*vsf����r扬hW����-ggix�s탉B9#�{�i��o|��1���-��LS0d��S� ��|��M���)>>~�g1٨�3�:�E�i>�E?=N�x��?4f�͈��㋓�9lV�G�5�P�~��3���E���_��v����šai���1�1}���P��>ע�-}�4w���R}���L�o��(/�S�����|�~�&����3TS �7Z6�@��()*�m��Oݽrѯ���ԣ�����C&�Ĭ_��*�����/�yzz�N�4C/�7�;b]���^_���l�B>qo��;m���De�w:pv?�Ӣ��[b)�y�oHz?��J���=/�V�W�:ǰıv���5Ԗ�C��a"]���Oވ��Q���{�W����w�fR����xs������b3#I�S˹��r	��F��Y�N��j���h�������gB��eGrֈD722Z,@��~�d�jt*���͑LVB��3�b�Ƃ�;�V��� �;�>���)[�;)�XL��o�Ee힡=��[a�V]�%���|��� /���,(��a���_󅃓�J�S>}�+m/����π��k�G_�e6��:�;}>���F��j��s���G)GYi��N#&6
>��{�<"8Į����15���>Y�WTW�%tQ����﴿oM2�-G}�_�Ʃ)��a:ݯL�%2�k{�7����8�����E����dQXg�K�W05��[c�w���S�^��91z">�/j��}��c}�*�������h\/�����>�i�.C��[f�P٩=��?�Jk
�	z]|r!�^I5.W���Z�k�=xBӱy���Ƃ����'R�������>��\��*piJ=,��1qL�o>͈d\�59�G���/SG��p���E�����RT��-��Ȯ��h�?毠h�<��eA��@f��#�����H��%ޢ&8ufo�ay=���%R� HJ��֧�"1���s�(Z�Ow�m�;�{���c)�>N�EGb�?*M�U����1�������+�sWxcb�&������	sƿ��:�m�V&rؐ(��vi��%G�����*�_���¯��&��Cg�>t5�D�R��;;/Cyeg���|�y��S[I3��}�7�Jک!Q�$�X�d�yi{�-�t�M$���+8�!�8�͎N���9��(&��<�k>��,'/oι��*�������䳝����:~Tj�q���<�cv�(2,QϚ�4�5X��M�wJ$Q���M�ԟ1av	'w0l97�æ��Q�~:S����M�+kn���ʧ�R��.���݀�C������ː݉9���0������B�w�[��c���N�_�I~�G'+�l��\��x�r�Ʋ��q�7��{���v�'<�bD��Au;-d�X�n�����7hv	��|_�DI��!F�*�m���T�g9�Q��/�fH ���\Ԩ�m��?����)�-�RW��(���fF}��%ٮH.�&ek�,rg�Of�Nwб�����m��}xC�gH��CR�i��:Y�f,�#�g�'m9��}�^�^P?�=�y*A0K?�5uys`N��
+����jj�0*~���z�Qޓ/�S5np%�ŋ�wJc���q��΁��:��.�ɭ���ԓ��I��!��n��'��ɯ����e�#�?�hs�M�i	����i|�����7o�ddd����@��u(Kڡ�Evj��Ǻ��m
��v��U���tΑs~h/h!�R�:S:5���;�q(����yn�J)Q������s>D��h��X⏬p~2ğg~�|�Ľ��:��i�||x[GGJ4v��d�|u�'���W�1o��xo���FS��ʬ�,�Ƶ���Ԓؓ7����n~���#���i���R=>�z�q���ki�H�������&��boRu�t�+�Ή�&�Y�{e?�m�*P��e����g�T�-�͛�X�L�G �%�;��4�U��].ڙ��YqyiQUs����ii���R��#AKa�X�m`M�$��럾�1<�l���~�ț��Ҁ�@�侕�G����Bl)�]�����-ڋEńɲMؽ:���n0J������S�7��z�%بp�GO�۵�+�%n�?Lic_t�Y��N�$�'l&72�.WǾ�N��K����zdK98b��7�M����t:A1ث�����'��]���B���#��v�W�p��ˇ���t���5Je's쵼���Uu)�\���!�S�D�i� ;O���$��7^T�j�4g���ϼ_��>C��30�6U7D�˾K[��Ȧ�i���1��*�6^��#���4L-���kl=J%�9�  �4>�Hr�R����_���H����Ew���~��	���O������w!:'��"���L�,���U��ɒ��K �$_W�?A�5A�Y�#W�(����$�S<��M�XT�� *���5�.�8�r,�$�p���(�K^9����WA~++Z2��B���tG�+ڻ�9ө��锫#aW����PS/UZ.�,�h���V������OU���Ay�	�P�m�&D��=%�uuw/E�Wt.[�d;,Z��b��9D�y�������V�=T�m�ŋ�[q0\(iJ*y��D���P�E�f��8_���b�vb#kv�v
�xbfױɭ�j�����B��NY��,�$ߠ�^{�]���	�U}�(���>���C^^ L��x��{M�%��ɑJ3��e%���������x}Z���0�O����d�Sbs�DJ_تʮ<YZJ�@I�ݚ�A���^�L�R�M����E~H�W�
�V4���=�	�I���jI��6�_N�_�=M�'�+��:���̣X	U�����
[ZZ��)���½����� ���
���p��Š�d
��r��u`+�M�-YDGM��[TI��ꢷ�0��{�h	+E�/��3�%&&������Dl�K�4�7�q~��̓%� x��P��4�Ou�b�.�
��R���G�<����cK�=�.\�&�>&@ƴ��e�c�za���U۸��aZ��p�@KFu\�vB���3_�׸�ǹ���^���_"����RN ����·���$Z'yˁ4a�����1޶�C�mBgp9�^������p��҄�p�'��+�/_&�X=I�Eos�t�v�%��
Um*
�𱾾�<N�w�ce�ؙ,�}n:����3꾙���P����>��\�U�-��o/ٽ��[q�a�!��<iQKj���#ݽ�G=XLt9%x��$5�ϭ�e��Mid���B������p�,��Q�2y�.Z���K�;!�傴�s�v�=��t\\�J"L��BVJ��N<6�꧀�ɲ�DP�
OTvqy���U�.�?g����7��fCm	��Y	���O��+S������2xD�w���Ic�=��_�\8,���԰Sk��.N�u`��5�[f��,o��Ud�f�Z��I	� �g�2ݙ��3���]�-�4�gw��u=��]k,f����&���n'�	��� s�K���8u�su�B���#����CCC4r���>0J���c9;=9n$��)X���V���hO��=2�"γ֙�޾Ђ���''��M�C� d��xkb�}�,ࠇ"�P��;��=?m�f 6r��MX�J�DlK��֭[y���{o��'ҰV��vn$�]��B#��(�6 sL�^V9��~�������f_1Ά��H�h�{T�_H���o��� �]�܀z�r�����n!���gJX��Ӛ���o)x3��B�e��E�!m�m��4ՁoC��ˊ�(+���@yE�'��ow��=<e��t����ȵ����t�+\��_<k�M`�x���c0lx4�������	`��=ǿ�����`�y��E�������e*2,|�B)��8��p��a�H�雼>����P�%a��]���J��o���ydX��RW���̍��A�����ν��F1�x7<hL	F�Rz���i�:�p��ҹ�9�pt�x�r�0rq�G�\�#,�,��۫�6��I��n/�z�C�da�;M���-�mSCF�5�N�M
���ےdj>�(/M����c�m��D2�@{�!���[��n����;��2P��T����?;��	�|�ˏ-�U�/�4q�t�S�c�ɧ9��-H��u��Ҽ���Gg�u�ۼB�đGU�<�GV���%����Q�n�By��+�,�,��
Q=���>ӕ��y@����s��^����OU��na�V�~�E�Uʖ}�T�UTL��<�Fn�`6��;hοG�|�à��.���1'`حr�~��߄X�Hĩ��n�M��z:+�7/T��6��q�a�{��#)��DU�AP6 u�.qJ0δf?f=��{EQ�2,v�un�,����������x<ӿd��!��c?&F�7�z�*,U�n`W����vѯ�}��"g7���y��,�����~�MbqQ�����F^�;m� ��������VC�F1�����xE��U{A�D�mh�t]�����V�������0�@TΡÙEX}�mY�J�cX�XA��(f�<$���{�gBdIKޠ%³Xȸ��e`����q�N#��ڎN�PWaV'�c��j�Dӯ
�3�;U�W��66@Ex������z��`��*������`H��%���uV��Ug,�:���~���!B$���e��E7��NN�F�� KX�O5��mG70�j[��4��d��A��F*�t�~�h��޳׉��|t�tl�m���^|�XL��:,fZ��\������6c
J�(�ՙ�x����d�B�ϴ��/9}��DAц�aJiQ?�㭞\�A��{�z(R��<E�ր���"���H>��u||<�����@���D�@w���ė���;:�`��DrQ>����_�����ax�"{X��t��!OW�>�%$���/�+7� ��u�sh�����2LQ ;Q.��o�th!�\�$��yE_ۍ���M'tx+���rh�z���)�M��F1�D@���6�k�f]bIAA�r:)�iT*��7P�����X�wߩ��-�|��P3T�r);u^��~SnQ8[Z�����]lq[H��<����<I��%����*Y��^AUxҗ�'�F��R҈���8��&���7�ܼ��7�%�]�:`�����b~DЅ����E�� Pp1z�[�].7�g��#�����l`���i���.)�l��<MJ���ćXg��������[�C��Y*AA����[����}�,i�Z���{�y��ԗ$L����,��h �6	�(�=|iȥ�F Ф�	�HA�~Ɍ�q��eґ�*u��~�����G���'��UB�>�;�Y	��B߄7��a�wSL����ms@�	<�<�<��-%�a����|J��(�5S��X�����hC�U���+e�z�&�=�*�8�PJ��=#EA7Ja�E�~Z�F�0	��x�����7�,�)���N�� n�<��w!���s���W��uuum�+��JΙ&sn��,b�n}I57�_�w4T[�.���C�,|���_�D�+wz�*��Ȝ��R�4:����W�X�� �/�oP����,�i3j��U�;�Uړ	/�=�+W�Jڱs?N�5Ɩ�Z�W�!��I���mD�Y%��,��f�PGL=%�P�oO$(x���m��ᑜ*���9��:��	su��)m�ſ\��i��L��5���� �,�@ �jO�xiq�+�5�;Ɛ�^�(u� ����-	�������(jh�M�C�!7�V<��I"\�r�������I}��z�v�������}d��cVA���|�(��^jb|��H���T�%D�VqeQt·4�|N_2--�N�d�-�'�$y�pF�ʞ��q�nEI)44�@�3�}�4��6|��ڟ�(�T��D橻�m,�4t�w\W��@�!(���b�\Bݣ�t�6��#�Ԕ�W�a��+�0�wa���\�1~Ok^-�}i������ݡ�O)����bE3�>����=��Tʷ�������l���#�[Щ���r�x���{���"*��+dF�}#b@�Q�'���9)GUBLtb���Γw��c�8�JP�$F%�|���PҞ^'4�;̓F�������~\��T���
����R:�?�ڤ���%>#O2,�殍�v���+O��5?�υyh	/��w�_�[�⡛����Ax���(j�@��lP�[X�;=Ĕ.J�n��P!��v9X�u��W���1dh:Ἔ�g�3�[a�u�	`]��_���4)L��3���l#��/��A�m.ɂٸ�P�ɋ��h$�m|�i�v� �Α_�8���0ZQØz��N�9��1������?�1�TX����g�B<ǌ9�Pͤy%�d:`d���C��g4F֖�]3��/;��|n4��z�׽Y~N�]�/�(9��N9a��ԪƁd\���'����kV���J��z���/�$߶�4��"�m��@w�Kt�C�5����Mt$�=�	�Q�edd,_�������6��Ww��T��y�4�� �%޺�k��ш�m�f3q�b5����0��� KЖ�ہ��=С2��GI�,�l���A�w�igl�����}�#�s�D��N��"�M��.�`=��7��x�
|'��S�^	��VF�(���L-�*��}���r$��dJ%�vz=�����b�LZR5�p.�
���E���$�}�����-��O�a�Y���i�,���gf/{.�{2��<J���������R��Q
m�o6����+rؠ���(R�a-����������|�D��nD!��4��j�|!�\y����$P4�ps�p7Z��)�weee؛Pȅ��N�>f�h��M)�vp��Xi>{?���K�^�X����>�]����'�*�o�n�\�AE���K�9�R9f��~�pbG��gj�ccc�}222;�S��R��7h�pv�W�l�`�z ��=�B��(a�:��u�����͵7	�Sk
37��&�!��0��H��۷�Y�t1J{�W!�����ڨ�D�LU_{;	�z.dv.7�ibB�hZ�͛7!����LE�:���E�J���4�[J��w�����5�pvw���4ɐ~�4�b�k���N0�jJHK�e�j�0O}���e��4t�-)���(�d�m���![���s�e��P�uj�Nk��f��A�\{fwO�����T��Ƙ� ?6�c��G<,?	�2���CA��>����]�QMG����"^��
笠n'��������s�v�kz�j�fbb�s��H}$6�h���]�w^|e*ԙF_&�x�W�?�m~R�x�e���!���)������Wmb�F+���b��a3R��=������썞���L�d�$a��M�5�H�pq�v��LvjB$���Z��+��vTVU�>ݝ��>*�f�F����G�),zZ�ѷy.����AkX)�������|�~1�]���ߜE�#�w�,El�i ��<UX�zr:c��M��=i��2�7��!�顫��6m�������3�vF�m��U��5�
������w�X�>�,��&9��t�z�Ӵ3rg����vBfM0!-��i���&����J;�ƆJ�ƅ��;`VЋ���?	ݙ��6��}G�s�F܏�U\94��Z?K}a:#W+��Pu��b�٧����F���A�	s;����XI"�J�,`+�q�PT�d#42��³�&ub¯�?O)]�a�{�Z.�C��T�{��pl�����4� ��z��/M
���~��
���|�ֻ��� �l�)��]�._�Ltwu�NTr�tr���?+a��o��KVR��bҼ�?�z)eO6���V��Z����൫���� ��&i�If��.��C����f\Ϊv�	-��,X��J��XrD��6_@�:�M4�D�/\J2=�����K�u��s����X�6
�����������@=݄�B+0P:�z�R5�pu��c)�s����ˉ��G�m��~f�Ni�v��#S��T�$�zL�6�� �U�7�dfMMM㚫����T�9��Wz�x2�)��]�����V@��%֢K� �ǀB�
���՝�K�ma�b%�}
&��s�0M朡n��| ��>}�777��V�Aq���&��Ǐ~�Y]�n�6�.����BQM��Ho�N��}	]l�@Y�]]��xY��5`N*�-�����e#�� u��A���`K����4v�K���F��*�����D��˂��g}���x��m��@ꈻ���E:�"�'a��S����$�y�8n���Bk�u��1�դg�?̫��%U�}r*��X�ø��Bu��F1!0*���3~c8c��A��=��>::����/qu��X��y:ő��O���? 09.�����<t�����gyB��G��>u����N��,�*�N���KT�g�3T-�g��������W��L&���=4D�}�.����S���0*�A�O����|Y�W��f�Y�C/s��AVEV]Q޺���-̜>)�J{�#��_'�:�uv�nnI��;�hc�����s�'����� M_Q��6G�����2�-"��S�oa�ܽ�'�xP��[]��@��9��W{��LI���&����b��3	���wї�O���۹O��ߝ�{U�R����:�sϰ �7~m�_��n�X���i&�}Qi��R����XD?���y] �g`q$������8�(�>�u��aŬ��F��+�}R��`̍�0Ѕ6O�����իG��*_T2P�S[0�� ��m����vM��g�N�ڗ�����5K�4���r�k�t���6�z ��_�JY���i�)pM���Bۑ�nV�y��e,O�������,�n#z��Dk,�.*��io��̓�'T ��Z�F\�Α�Y��}A���?��5�g�����G���>&?�/y��{I�nC_K�C���m� ��wyys�����@oqIl%Y��'�I,H�w�9V�∪�O�^����\�}���G���t�0��)(�6`o�Em��Y�f����Nx�����4D���
�!�|��F{/*�[A`��+�#
}&��o8�?Ν��܆v;�ura����j C(�1�K�$�$�UzF�7���HF�0�(5�-�%فn4fz�mR��v����C!A��m����`��+�Ϟp'�Jt��
�d�ީ��?�����6
��l��Qj~�'�'�u�>�9��i7��O~-[X|�:b���Lz����7Bm}�J[uu�#�vB�0`��ގm."<A�����E��^��S=N�ߜ�I�fY�$�h�Vb|������j�q�|D������W�&��7��C���U�xX �m���Z�R�q���ŋs���F �o��@g������͍�>\�D|̳�r�v I���/ҷ��h�V�D&��'�B��:>!��G�|��͓�<Y������$'����5p8_�<�Rˁ*Y�lr���©N����^�wd���(�^NoQ�F�$PR"�ϡ_fwk�D>���{������K2G�D�IT/��sh���4D��H9��+/�JH�����"?��Qz��K�fD�1�u��2�����ӸCLN?��{��l�-\� �UʧqvϞ���# �觷���{R�+��_*x{�D9���DnyL ��Y	�\�Л���ԁI,e"�<}�D�����3�����}�=;ru|az`2.)ieapp�=���V蔿=W7��#}��r��h��&�������m����x!���d�&i��&���L��+-��A�O�-�\d�P�-):_x�J��͗�yw,ŕ111���,��d��]/�_���l�#dfe��(���/\�7w�B�=��8(*�I�5�4v-�F�%���#�w�z�ҿ���C�SP�����Ϧ�U���hsb�az��@%��H��Q��Ѷ�"�Zn*r�-��3���n�L�?-v�
��˟��5ꩃrBF����T�����Ν���ݥ�&�w�z#���^�`��2I �n{����ϧ��3�j��Ͱċ�A��K�ɿ��"wZW���!�>�vӌ��p�힁���������뎔�9Ӗ��n��?
*"�.���Ǐ�f�<�����Sq��8X#|K۔)V|47IK�����"�������ù��I���ߊ���<��5b����}��]O�^��QefɊ�ܦ7��,��=b�.�X}�������ɅYi�٫^�r#��H���	�8�jS�!��+!��`m�ddP�mQ��v���{���%'#��ΌI�b�qJy�����׆�}�D?G��n�hf.qu+�W�3���O�<㪢���aޗI ��ɛAk��Uk�a�n��F�x�r��M����? ��,��Lꫣ �b�}rOL��5Ð�aX\oO�G߂N��"��>Y�/�P ��=޴��CZ���xkp1�D,8U=�FR_��������
k�ۯy���¶ˢ�m,^��R������b�>���cy>�얤�=�\Ǯ�r^u���!�I��<]㟐��A�^���;\B�1���rz_SS�ι�%mܾ�	t{[P���gL.�M9��{_dK9g?K��VZ�`w��T�'�,��Va3�' `���龳�Ȉ������y������2rAW��氉H�ݗ6�L�y�>�|�KDF\삤9�nZά��r�roc3� ⋳�aaa7�a�M���"���ߘ9��,��"�;�)����%-O�hmm-IK�@�~VD���$��R8��d�d���3���勝o���"������dB
 �2w�n�6�]�*��@i���_�~9�>}^B��$on�i� Ž�xqVr��+���s����a����!����W���1V/�R��P��)o��s�\IC:��΄\��9�<@���:)4㱕Q�]��i}}R��.wff��"�,8ωv\>4������,�E�i�R�_�,���f~�a@2@�!jsW�VM��C��b	Zr�ut�A���FJ���C�<��B��
�.����ǫi7�۾y9 o��� Tzc��H���Оu*�_������$f�ȩK� ���?@7��>98�Y�6"|�4���
��zn���2�}��YȰ� �f.d�Οkՠ��vy+�>�+�]l#o�F	�
axh��C�Vs�q<��S�F́�.���杌qF+:v�A�jb��4�A����-Dٴ�i$ͧ�P[�D���������g�ك�7�}���J�W��D���jލ���-vsy!9���B��mSoN�!��|�,�~l��ɋ�XEH���ȇ�牙��Q�ǋpmZr0'''����&�+U2��99����O*����m��� K�۝�o7�x;r �����6��ɽB�/8����C���-\J��S&h��(�4uww����(A�y���t�ģ	����)����u���(�"�5�����2�0�zrкw��ŒL�_(C��x�FB�PK�ܹ�Z�����5Q<���T!!!&ox���T��ȃ���s�{�Gq��l,
S���M(�m���%j�ح���Z�oC�Ȣ��'+[�q��L$T�|D� �§�f?��+�)�S�y��Oz���P��rA��g0k����#����g�t���;@�	r��p����ae�I�*��r���
F[*��\G��Oޑ�(2��~ �~?nY��X�AQՓ�����ŴJ�Ae3��\Csss?xhߐ�2Kz�Ei���H��翧������m� �7�X�n�Þ��YK ?*���#�/��.���$*1��Dn�a�	���!�Y�2Ɨ�hJ���(EZ��夰9ҹd0@���c8� �=�Ʉ_�������L ���<99� � �1�m���S3o [�ڈ��y
)w�i4�;A�����y���E���7hIjc4�����B�����u�>��4��a�7�0�Rے_ul2��
����Ͻr��O0�tv~C]��iL�9�p��d��=� |ҎCn�z����ʯ�Ku{	����3ݗ� ݟ/�XU�B�'���n��� U�p��*�]A{�@ݦ��Β�1ǏW��7,`vl1��m�a���S��������f�<�9]}}"H�KLӟ��%�AD<@��҂�e�S����/��w2�?�>q�l�hmm�U?xpV�`�lA�-�
�>��A�}[��ks��-�%�f^�"[����}|����,�d��db��5���Q�"���9�qh�h>'�����7�l��0�yW�M�8=�ʀ����%��q�prDW�%�c�"GV��n�az^�S>c$$$�c-�V4�??E�����ʊ
����J���c �����!}�⹕O�e��=��J�������P�����Ǚe=��_�~��®M�L��~�������`�}�g�!�2G��5�����{�w@�y9:RLѓ�g1�xaD̛@���M�KHH������4������;�|��ۡ|�vd�y�d\h������.�Ԫk��R<� ��A���([�+�f��0餴����w�n0}���K}��<)����)��ME�����{u~%�0�ߴߡ'�=!��e��U���N@o�A��ӷ�Y��
@z �5�M�� Pe|C7��I���D��YB�gqi��{����?K���_ ��C����?��a���0��`�sD�6���I<��F�d�"�ws�����G��>�X����0:���1�芆��6�j��;"��sc��pG�W]��:I��$����<߼LB�m6S` R 
�yϦu����N~]+��J�C4�bv�]�ߎ
��`4x_���%J�4��r��=�����z�Vj�J��"��ʕ��j7 ��=�!��R�}�'����U��y�pqӨ����4���w�0������+�� 1(en(ʙ[�� L�N����z�u1D���w2��n{��*��C�.��a� #����NrH�i,��>�`�2�P���|5�z����K��ECt%�"���9^а�Q̡�������� �"C�����`5�0�9��I��X=$H�yD뚑h�K�M����X���0@%luu����5��C�$��N��=�ʛYWEs��.<�� f3 r�h%�:"��0d�yu~���̪�_@sh��_*�B�������I�!�ܞ�ۃ�<�V����.�C�#ȗ/]Z���}���蝍�"œ3��I��!�쉾ïE�����m�0�P@1��g���<rd�=��c�p���{��+4��K�ݶ*m�'it� 7P�$z�!����L��x����Ƚ�_ׇD���Wٰ*� aZ�O�VeC��˪&0���Z!9��[J�i]]�\`V`V��iG�z�U�ly'S��>�G��I�(��L~Q�^BQ��K.�r�:���B�����M."k�XzK�'-}�b<5t�{��vUt��d~r[�V#mo�_uQV�AJ�bs� �n� ����9HEY�����m�>7��I��.�X��~r��b�������C�9q=g�Tx�n�[�������W瘚!�$Bڜ=���o�B�R�`!� t��s!��Ͻ �΀��2�'�h	�F�Ɓ�MK�âEi��>ri�i�i��3�J.�y��t,M---E2��8�/ �'����xe�Q�z~�.<�
3J��b��P�4l7��jʊ���_��g�o�v��\}kNT\
�JeT{�rM���/m*�TY�o��s� ��@C�P����bt�5��|LXE�
s�e��o90�&��!�H�.�/�\Ho!Ĝ���J��d�rP�467g�;%W���&�Z�X�b�2߼�{g�^�N8��激��[~�NLL6�;�~��Om�'��0�}�^X1˾�p{CQ�Un����m�D����/��?����}}=������6E�Z�@���*@����8�u����TQE!SȈ�O��Ulz*��͍Oo�ܽi]?>@]��]3RD_��pォ)�=V�����pߗ���)W��gmh�Ԩ]u�1wU{�.��T�J�"�P��N�"�Ko)#��(�.~l`��� � %(F$��j�(���h��ס���������9����d�O*�8�D��O��Q	�c�{�����lyPܨ�oU��[�^�Ԭ,27��,��<�w��.Y�dRhb��(u��"6ɻ�%�\��@���K3 �Z��R��SN��q�+�{$'�.k�
�\^�{y����	���:޷�	H�e�rL;��D��3z���N�����x�6�< ß>�6,n�p�ܞ���3288H�%���;Y���I1��r9d�Cz��}�:p~�\Ԓ�5,��
�Ld�	�0%�R��a���9����R_PN{��_0F��U�U�	�jܗ�&|��z�pܳ8��P/u��_��� <Odj�����'%$�5� ���kU�șq{�&���ͱ)��7\�}�p��I� �h���k���P���? �0�U�����}�re�Fa�[�����Ew��Ukp��y�:��0ԯ=3����	�*c;PY@��&d/b�P�/�*/Z@{�?m�Gϟi�;p^ ����0�7����_���-r�k>��Y�u�Kj�Փ��+@�~����C��WZZV�1٘)���G���谂�b<FCbՋ�fEI���C�:�� JM��	�'���w��ע	oG7�K8 &R��*-Q/������1��A�dNI��A`n�o�I����"�.�G��Q���b&�l�=NM?��������>7�:�Z�����l���.rB�[��Cb�P#���#�؎�w�$Ԑ]�J&y��B�ʔo[�u���2�_�+	�W�����~�CcH"��}
/[F�����3ZW̲hT���c��!	L������Χ�8����R�����t�ӎ;v��1�RD?� �r�Sl�����8��x�9�����tP�M�>B���� ����I̒��5���8�[F��`Β�S ;�ZUy�������r�D�ߩ����:)�NxE]�8�ɃB��ݟD����-�����<f��
�ʚ
�#��&�e�8��#�?=q����&���4H�'m4�)Ed�O�gNG	�>%��ٿ@D����Iּ����Q��d<����v�c���E�c���i���ifY?f�C���9XE6�o�R2�Ѩn�M;��s����Y��� )0���=#��9�ʓ�pcS�h-<HgY_o�FU/�A�4�u��i ��w�O�@�5Q<I�vy��0C�2�H���<�g�XL���ܚ<��p��$��m��t�d��u�6��3(&�]�̑	w����Y����b&_��Peؗ�=�Jo��)--�y�����H�Ul�vh�3;��:`��N�|�g�r*g��T��
Ӿ���L* �8'J�O�8[�B�E��
0�� ���N�P!m����
���W"?��D�0�H5)2���@��f�q��О|�nG�D��������$>ޗa��C�\�b�ъ)��0����~�_dmd���D{��cR��^=�D����#�&�����p�[��Ź�� ?�B�`П�����lϣ����]h3@p# ,�sss�����jS��*p
��v�H�ʂ�S�{J������$�Bg�	��1'g�I�3Ψ�%�78�˖�����f."���A8Zan~�z��z��z��Ja0��m�X��џ��^#���}�%�3�Dw���6	���+��m�=Q�q!�(#�S1�}����>>��d��7��l.}>�諸�њ�&�d6V_!�;�P(Scِ��mݐT�4S3�������t��d�B�܈�#�c~�f瀀 "����@���>3���/-*�z���w�_��۳�c:��mr ��)!�lV�����W���F_%$Y��D-��/���t�gE(������{�7�j���ї��������x����)&�U�����1L?|���Q�Q#�2}��ɞ�UvcO��	���{���Ԃ�{Ԣ�����(]���O9Z��=�ɻ ���W�?�ȉ������6�v�ax>i��Z)xQ���0�,없u��G���|J#�:ט�c:�|�ͦ"Uc���ۨ��}���ڙaSy;m�K"3��|@�0/S�.Ϯ��Y������<�V�뗻�f��	L�0�M������L'OG���I\�B!�VFB��a��@ʛ�f㯎�'�߿_�6��x�x�5�&/OX_ut�?�yXSW�6�>�ѶZ1N`E�`�8�d��`�BFdF� �<���jD�(ATh�Id�bEP�� �2
bd����ɉ�~���w��{�?��pv�^ý���>�lQ�i��$��~�a�H�H�r�j�N��$�9,$�D���ɾř����w׬F+o��G�����[3���4{��{�:v`s�Q$z�������f��#m3��I���Źs(J��KJvμ5��;:�����{�!�
�=�I����M�՚���x��Q����m��h��hkp���a���n �peP?�Z���sYYY�.m;?��T��q��b�����;7�����ώ���vF[�8�����:��$���U�
r�9dM����EF�������{�J��/�r�}s:&6��ь��qX�3r��uK_�h�������5=9Z>L8��Ȭ�cT�Dw2����h��������ӗ�]��ëK������;�����6�L}���mY���v������S�no���ǟ�M2L�An�&
���D��dXv�Pk��б��.-��uK�;���ۓ��[6�Q�qͿ��59��a�"xpNN~zT8	~�)�i��U��>CCL'!��G']'���>F�H������/b��}�	��e�͞�7n,M�i�!���j�	(���:��>X.Y<3��a�Q$��R衼������5:�h�ɥ�w�����9��]{�z"���CC��?�ŋ�#e���n��_� �I��X''��߲*ͷ��M�4�����������zFڡbt��-��ԸH���vf�?r��DRg�_O�k�g�#K��	�5Z��_�6�VuY��]n��w�{]��Gl�EEER)���xzg����5q<`�U�SN��4�dt�;����ӟ��6]+7�
��w�\[� �<�xxF��ٻu�ɓ'��#I��L	щ���!~ꭂ�\;/95T�����O~���37�X�"��4吴�����������"���m�K�������OY�����{/�Ժ�^g?*v��p�xy{��Mpy��7gd#����]�hv.,k(�gӹ��Ш�wlP�������'b�R�A���z,�-mw�1�A�{tt��q��=vd��JIh����X^����Hc��c&�T>�5��tS�鳛�|�'�Z� �����\�G�%4لϤ�!���@�{�����8��;�Ҭ�bC�R�$�����-���m�Z(Zy�<^�% 83~�AG���˹�Qf���_|?��l5^a�� }�oJ,��M�$r �7Z}�;9m9��7]�mX6R���9�b&s�a�o�%PQh5y�[�g�H�UG�&�%�C�k|@Q�P��}�j�������};/o��\���^��rG�g��z���(�9"#�V���Z�Mo�y��<���J�m��I��+��2h�h.��f'<�O�>o/�\J�m�D�I�?W�?Z�R��ۺ��U�!�A�./�K{%B�9��æ��(��BÊ� ��_��c&��v>�-��S�jQ�~z��uѕg�`��7`�������Ѳ%�D�� ]�t5�<��L �Ti�2̵ٍ32[��<�#������$�oqm�'�ϫ�Ҫ�P��bmH͕k8�R�S������]�頻��hY�h���ݔ�h�4��"E��q���Z���4/M��`ck� �ޅ���+w��-���L�9���Pv����?��"��뫆jk�e�k�~�GHww��//6D�%Llv*��ah���T	R��� �2%�������!���Y��[e.��^��|
nG9ѿ�H�_�B��N�-B����JhKS���gF�"�ۗH���ۺ5��z�����(�N=����l�x���䌄,hBY��c�":����j���ڮR�d��u�Qc�?�Єb����c?i]���ѹ�����s�g\���Pդ���9 8WS�9��'T���EE)x�?M��z(w�8�edݒ�HT_��4�A��b�n�����,�Ԗ�R���2 ?�+6$X�!`�C���@Q�:���!���w�(��� ���bQE��S�Uo�����.��u�w�A�/��;�F��62ԼLLb�UI�=j>��>Jrrȝ*�F(��j떟�b�y�4Լ��uQ��1o��5J2x��=��Z���J�-Gx1����L7k��k�������D!R]*�9���T�}��C�^�z�<��5ڻC!mbr��PT+��&���\�j��W��n�dZ�v���ˢ��~�(�E�n/)��yad�*���O.i��GC�TԆ��4�Ri�66wՅZ�,���u��=��ak�6Q���@�//��x�Sߜ���*v+��l���ބ�U�W�r�y2>�����/؂ |�?R��a�O6T*�^{VZ�c@s}����j�,�e�)�SPL��������y�L���E
豐�L ޑ\��[e���l�s(uV��=�Ǯ�,]�D�_��PTO�O�����Fw�B��(�
J���Bd�&����P�B9[[ۛ���A�N' 8X�İJՕU�[G����1�r��6��� ��JPX�j�VDC���@�B�9DX�I&''"w�6K�;wN�Mk���2RT�K�p ���䴹��^ͯE��/_�loȰ41v}��A.�&��$-A��:�읃��ӊw��6M���qAY_6P�O���$l��[#���ޕ���,���}|r����uW�=�yEɶ'ߥNl�8�w��Z�w�3��4=o�_����d�o2ɾ5"�e�a��j�g'�&�wn�l~2�>d΍م#=��#,���l$�ܚ�V�Ҡ�U�� c=�N[�p�Q;;���_`�H�:�MQ|��FG;��+�����L���쌹zu1BO�Ug���m�L�:�3H��Ϡ`��_~izzzl���0�:N]R6x��W^Z�U�����2��<�����Qs�w�����Q�|P�q�{�lJJ��P�l����ڊే��;+���w�����؄�| �=��,|�4A�mv8��~��{4��~�j�R���nn?�>s&a]���7��^��D2D����_0���"����7�L��H��B�s�Zą��9P��'���:���J ej=�q���ڳ+U�8'�������㯡ms��,h>�=6#/oEee����t�t��� ��;Y�����	�)����ޘ����ϟ߮;xJ��H���ciAAAFF5ǩ9���J��g����ʃ�"s�Mq�*pt�CCCȈ�N��W�7b2��+�0����X�9E(G��Oc���X&Ky ���� 7��ۗ�0���A��P�����/P� ���5���D�yc���p櫰j��y�P�)@�]�����A)���T
%�.��447�CU^�b��_�j�-��a=��Z&��
����a�4��sؖ�=0�
i�~Nc�m�
33��:c�GP��s_�j�	1$���������ROf���L�vV\V��3��,ok���b,|�~�h0ǅ����ٖ��j�=�H#*:���w��TKZ��>CU*6"�m��2 #��WSm���jpj�k��� ��&�m����^�EO��˄�1�o�y�ˏeeeG]\�Bo��3L�x�@�����PM���:8;���U�˹�G�BQgQV�lls�ȏ"w͝�񿔶:���}}e	�����B�Ag'v��.4e�%A��V%An�/�� �'&%������B
_q=w���>t�6'On;+�=��wGf����?�t��`����|��/�����f��c���3Щ���w�?�JQ�����oٲ�����Q���~MY-g�p�
�S4;�P2`�S���������>/���%%��Q|���n�"�svV��
��
ԅ�#7 �S�Y5zcc���_<��h��!���d.;s挫��"��B�+#����XQc~��֊p��������h�u�sԽ7��}l�ԍp�546�C��
Z�E�LmEQ\��.������R&��i�� ��+W�B�K��C轍��4
��eF�g\=O�w�ȅ��)��^�q(M��CyCP67���!,��{�"˜�U�6�=�G��]�_�����@X�:4��!6`��Wv���54���'��d�fdli���>�|�9�1#'G266�j�����q�q�"����z�C�r�޾+o蜤bY{�Q��k���i����=������#(���Z&!���|��ڈ�2�J ��xj�ʕ+�����]S�TJ������.\� %-��x%i�v 0����G5gfFK���Eb�ő<0�����I
$�/G�� ^[vɒ%[���P�<S�����ii���$CD	(��e�z
>������i�p����88l<}��Qk�c)SrPWI�Z���2�2����i����K�Z�9��ޖ�u�9%ӎh�*�]x4 @ыe��IT���ǐѡÕ��уy��wzM%���99��2x�5x����"��e�%��*��+��F�x+pY�`�%A���������ֶ��ు#���{F&�	�&��I�?}�P,_�rM]vժpD�P��Q P2.�}�d�UH<�DoDDԍz	�Y�cЮ�x{�v�0��-	��NP���B1���%3��I���nY4/D��[�PB�c`@	K���C��P��"N�-~H1.�+Fz&+͋Ԗ/_�ޔ玲���<�s��i���)���wRS'��ii�tx_�b�����s,c��*�j��x���[�n]���Q����ɧ#���{	�Z��`�rd"�Rh�j���u����|����!Zr����_=��s�2��			��R�ԉ����@4LfѢ�`�%�^*�X�W�J�[����yn?����om���)'��bhz�
Z�1��O�b+O�I��j�h��I�i�B*A�EC#`1��D������zFn�v�4k��g��x8�<���x����zFo�Q���uy������ݻ�'N���׷9~|`�S����Le�0�PD N��X*�A��-��1�Wo �@��E/w��M"���K���

������	���~E�|�_}AQ���!�kc1n�(vxG���d�[W�jkˢ�J�٭����<Ӕ�&�uz�nގ>f�����`���_�A@N���e��**o��P��\K�$mG@f��Z�������1m�O����ً��j�]�^�&��q[��K�-�Qύ�=��Fb���&��ޫ@���+{�����F��1әj���rI!��ޔ�1�������-}�wo�B�=iZ��Wz>?i��]u���T{p��cG(��,SD��z�� zN�`���%p�P�B����a�Yש1�x��o�*c���dZh;C����MN�l�ܹ��nZ.�Mٸw��3c� �y��}���f��+��q`2G�ׅ�$�����>����p����
�������!V�_�xQ�_Z2#��>���1��eY-}4O���YV��u��8�*�n��3��b�^6;�,��XҸ�}u�����L���$����3�OK�q������Z�	SN�Kj��͌:X!�]?���r�-�B��,�<w3fS��{+o�;&�z���P�K��d�;kr��S-�̭�{h�\�K�vKz�Wʡɒ�kb-�nh-�ܹs��ڛT���x�%�D ����k�\��bQ�Eu��ES���:f�৫�����n����#�[��M`��m3���Q��VP#��ɼ����f����8�\ӑH�����@���n��!`b���������4���ETg�R�x�<�{��F�v�?�2�h�U�۸{]���t�����/�t<��,�^3�Y�7�0^���x�k�FV)u'���}ҳE��mv� ���{@Z�t���:��4%�X����Co�@/��B�{,z3f�{���L�NF���>�&��m��]�Zp�������AE�c�����$�x�4�����<�kXE��·C̺}�^�RhnԩK�'uܕ�����l���3��?��(Ċ	�f��u5�	��)��]�:�b������
�&hU���,٘��<�Ӆ~'���b��xF�&���"�fb"�ewo�i���on��'k-[��?.Z.��1�>�:�����q`i�!;v�N}�!����k �86����~{����̺��r*����Afݎ�u���EW�\)Ki!�l|���!J�˜�q���~�;$Kzf2Ug˧��\7׈>�:��^S*����M��j�w��JX��� Y���ؘ��ð?����+�$(���v(��g�+B��z�����_.~���○_.~���○�]�l��<�p_.~�����&ǂ?�ƿ
�W��X!�|xQ�W�/��|���˧/��|���˧/��|���˧/��|���˧/��|���SHCސB�`����ݹz��&��w>^��|�-��Wت��N�Ν�=j�V��),�n)��9�t����[�Q�ϩ]_��8,����_5^��=f�M·֡?�^�ݓ�7�v^��r{���oߢ�?Gӄ�����(�{��z�T���/���R�������������I��'� � U�`ݶ�������~�杰�q3���Ʒ�j��g.�Ő���l[��қ�|��!��C]]y�=<F��7�B����B��/�吪*-��"�������$� %i��6������|��-�I��4G��-=�Iڈ�
wʙ{����.O�r:h��9>M� R,�v7Au!���?�e�#𦯵�翺yY�u����?ۺ˫@Qd�σ3tBΘ�>�����_��i{9�&�9�r�5�\^�Q;Z�h��[��:�">��*��C�^R&!+�f@}�E�9B��ϒ����I4�������?��������:�
݁�E����'Hy]Z�uNQ"HqK�O��W����"%�u�h.k>y�Mj�x���;����3;�7���M��`��{��k�T��!��- ��uujτ/!�C�XdZ�<~�vH�=kw	|��E[|��/��Z<�R����b�H�tCbӝ}��1SwA^?���g�l�ӄ�gE���t�]K���N��ލ�ݻW{�*4�_�������~�������^x5��a��b���K�#��FdL3j����N|�w�p��0���z沃������m��y�{M��~b��9�*El]�g v�	|�׊����\O~�.1��S�ߩ	��|��*M�b�M�ޞ]�0#���g1���?44$q۶���z�q�֭[�%`Q��V��
���G���bQ�
�ñg����1RNJJJZ-ŏp�K����!c�I�8%�ڮ��������Еb�|!��^'ш���>48�c����9$���v�Fm����J��w@S|��������鯲����	FEPq1�3(��7e�`M_�6���}�����}�}���>�z�����LjP��hA����2��{Q`��SRS���K7p���job%^Y*��Ou��Q;����o��W/�W�z���c���G�R��Əa�6]A
]��@���+��Ж'� �d6_b�B��8��%��8v옾���(D���]�Y�`36�M��MॶLd��+��wy=+@֖��������sZ%�.��Q���Y�����?�< kS&�!A1sI��7?����mXPI�~&�N�6���_"�'���W��%d�$b�Ow�2�ד�َV�q�*=��p48*������~s� B�["8Z[LL�X�P�����T�kE�I�XZ��K�]��v,P�i�Xd���jv�M_�M._.)��X�^�2#�4h�#.9��z�*�e�_��0��/��E��i}�T���^#�:�ho�X��o��Q|�l�+,�z�C2�WQ����h�~T�q���®��~�:���]��,�M�{/���e;��,�w>|�LصClW��`�0�"96��S_UD�� N�ӂ������Z!�j8 #d��-��8���?�ˏ?ϼ2w�+Ne�֡��TH��h�`�Ka�cc�5�� ^�6y���嫒�nv�B���<wx��Ŭ��\�������-v�;�z���d�.YH6璂a�&�E$�+��w����rW�q�L��ܷ����h�u��2,,��F�Ɠ�s"���k���֑f�M�Y�#1�~�Yݿ�aI�y��n��z����Qm���7�8��p�ޝ
���!z�$�˖&t8!ҡ�v�BJȷَ�g	�m�F{X�
�������m$���ߞw��7~JJ�$�����V2�uw8C��lֻ8&��b���"��CNt���.fu��YU[{�<��������s{웝F��x�ʑAud:�]�(�:�����s9�S�A��%�1x+��ա�x���'�O��u���Ѻ�+:��.\�c�Ĉ�����K�E�:���"���M�w8	�K����L����#�1BH^FC�`��fvcoK.��3B�ޣ"�$���C��������I�C��t���zp�������zSzvI������!GHQ��*����ڔͰlV��%r��*Q����j̠�#�L�r�e*�1O�1OԢ�5�a�U{d���D�\pNd��C��H�+N��9�Yw����"u��	CJ�ur�ѫ�n��B���.{�'����l�(�V���G�p8J��L����c��dait�v]��?ڧ��� >Ml?y��l����v���-�و>�	�NK���Q3f�>b�C�r�`)м6��1=���	��;����K	o���n#}��ź�:m:m��v8;4z�kK�����%}��>��e':6/�������`�DO�B����-L�R8H��k�86D6�jұQK���<)�� ��n�e��M��^�J�������O~�z�c�Q%h܀��W�S�=C�*ۻ��߈>�	�:�&Կ�Ʀ����w�L����V(�L���̞w'bR�%����]0�ӧO7E[x�J�i�.��}ߜ��[��!�߂c���D�s�%���7u��i����(i�ouy��x�X.(����ˣ5�/;�J&���ry���l�qn"��`���5�'�㝰#��Jƻu~s���{_��z�Y�e�LD9Si����Lv�
���W�%��aH֐$�_\}NCz���߰&������հF���N�@��YE��ty$�ꋲK��
�_Z�����nXD�8���M�t S�}��F/5���i<t���*��Y�?L&�6:F)�|�� ؼ��(�� .�t�K 9剚���Oq&��#��"i0�cD�B	,�%*�~s(^6�����6A�)��m��s�<��	Y�����:���)����q�����v �x:m$��$����6�1��<�A'�_�|��ZK~��i�v��R�\UB4�kI������ۍ	��{Ж��9���gn�sA]��-Mٽ�7	����No^�-0�qƏI�KZ�F��
�ۇ�ޢ��Ĳ۳/O��;�&͝i}��S��3駺k��/�*(�<4���P�Zɹy3L��+���0�޺mυ��9����|��,Nյ��3���i�0����4�Y����w�%M�u�1*R�0�0��Ǣ�޽{���!�$Ϝ��@-��nt��I��؊�FJB<¿�h4�ƭC�5N�k.H������	�������b%��ܸrc&�&�q24��� �
s!9fC�s��*��j;4��i��@�����ʊ\���9*�Y
qt��F��%	CJ���N-]���,YB�S��r&��5���ڗ/_jeܿ?����}2���i��I0��������$���4B�yA[��w��p���':ke�\�޼~�>��.��MB��� ű��w3��R+"j�/�{31���{@ӓ��
\3y%��	}�w��j��h'W��+��PN>z�H�`�-"~���?q�]�����w�z��j�"�d��znTpc�8Z��;��L��+�$;cL��ǯAk���H,I6lG�i�C"&�PW�����]	ۯAF��_wx'�q� ���d��j�B�)�eA�h�tZ�d38��Qq#۱�n���4�i���N2�]�Z�}��'�y<A��C8�0=�.�嫞�Ç���Kn�p��F�Q�6?A������Jr����v�~���@��l%n�TE��Ũ�G$�=(�v�CMM�/� |k�E�}|wӻz�L�gR�S�EV${��1�Nл��r~��K�����_ze��ݗi�,dƍ��l�k�	�ȝ����)��i�?@h��4Ӹ��'y�v��MM��ٙ��S�d	h����c���i]���j�ˉ�������A^NɢԘmD���(���D��EZ����>�����X��8�*�ᑀ��ޕ�[i��\v,���`~�~���.����/Bͅ�cmE�QK��Zl��`r�[��5��g?61*��Ba�Yl� 2��<6�ei_g����V˸~d��H���}drz�;�e���G;��&!�<R�{P�y��<��.ȼ��p���N��{Z�d��R�D�(��z�ѻ�f;��poL��G�+���Aiw��Uvo D�R��2&��!L�S[ѓ��p���J*��ǜyZ����urZ]�n!Z̏�d~!�}3�ۊ6���P�-nVb�H��^�`P���FR������ׯW���!�$"��Y+Jۮ��z�����Bi?�=�3}hk٨c��UG;�1�7�2����C��i,�K�» !��!Ӹ�l��&�V�&���T�"����nU�֊rɾ8'�/���9�p�I�yML�삤�tٍ����X\��]y���C� .//��[8���3�Z �4F�DY�29�˨@��R���~�/�v��B$r�Fj％�c{�]{�5���!��0�ג��Mh�&�D���3SLk� ���F�7�3��P�W������8y;O�������n''m62��Ԟh��=�)�Iu�cED���꯳�
��c	��IS������,�U����f|�v�l�;�XG'r>���F�VT-��Y�Cm�J+`����x�G���Zx��x�Q�AsFz�@���H�}��˞,�Xkd6��D���y�E���*�ԑ�'j���J����&��hn�BJX�.�	0RO��M*���uE�i��P�g�:le=r�u�#�ni'g(�1;ژ�Y�~f	bE×�V455=a����N:�Xi���Y�=��pʐPft0333s,���v")�v��iUU�>�r��.[=~amz��tAἁ��Fe��3
Q�F����Y}�t��3�qsP|���k߲֝����c9��}�iWd�qW܋��>ZDV�g�쪯e�k~B;�+�c���d^V	����G;�ʙY��		_��W���Y`d��M��T��T�����*KX�Q��w�3=m�;���.�޼iS�$��Q��mȝg����p�B���r�8��t�A�I�.[(�1��.�GFp�1�3F�o�o��y�����WL[_<V��ڳ�CJu'ù�8-��"�I���p**&�PP�[@Z݈�d�� ��o�?N�z����{�ky�w\����'jV���L.�xد�=�32S�/d���!�#�]�챀�~�ظߡ��"��!#$���%��g�<������hoIl���������+�&�;tZ`aj�&�*}9��N�N��	Z����	Ov�1�I��7^�k�
�Wډ�h�z�wb���n'�˝��^�tZ\�-�^_%����+��r�$����%�����(����v��/�Z��!X����	�r�Q'�*����ۈ,K��_b���d�]����F����lR?R����1e��7]Y��:4�ot��co%|s����<
C��$��܂ſm��������|������B�8����,徖:�煝����������ӃA�p������D�S|�;�D|eψdapSk��I�ȝ:���:M���c��]qP�����	A(�⸲i�@(��s��L�;���ߦ#2D�zڻD'��M��ˮ�y`��{c�Wճ��z�
���(2%S��Jl{g�kE��O��E�+:<��aKC��U��0�l0y�`��y��p�Dfuͽ���s$O�Z��)}�Ԟ:择�\���i�KǇo��0�hTDB}ϴ��9V�������IE��AD�!K�g�j�@�£�r��$�!����cI�|�#NP.�����~��,^)W���̠%r[�[ᔾyx&x�\�Fx-Ӌ�g"�B�ĊZg��v��/<5O��RT����
g��)؋���N��V��0m3L�?����9��:�k����J��~�t��r3w!@w~%�e��x�]1*H<��bv��9��~�o�����q�1N�] �2ΐ�^p�ҟ%����Uuj(�B�DCI:���wF�=��}ѽ�V�*�;_+������?~��-�D~_��_r��޶�♈ C����ُ�5k/��&#�����C��a3vװ(���އ�^�Ȳ���D����)$�y�N=�c��"��cG\k8k�X�\�&�B��K��Ђg�-��c���r��~�K��J<S�g���:Q��Rsz9C�W��SO�#�N-&`y����OD��X��U����e��C��.�)ii��u��Q�^`��<����a��dB���뙰r(�e�C��h.++C�ύ$��4K�u�L�]��vE�!�4gtr:M��]<�mC���bj�%R�s�����8Y�Z����!6����O��q.6޳<�gb:��l�V�2�Lf?�U�<+�����V�q��w碚Nʐ�6j�Xc�x�� -����;LLG�D�{U89�&g�����c�N4�VTT<$"�Rd땐˼uK{��i�s�����a,�yJ��N(��Qv��2-Ea���j�i"�2r{��T�r�RĢRf��z*�:�1�y�!2d֡)@����U�ȼ;M����\�/�
��R�F��0w�[��U<ގ��33�������*�.��bټ�5?��x}��d�!~��=����ZȐUnР�J@����CD�+6G���n�͗N9V��ޗ�1�$�Y�`�U�8�x����gW�Yb����B��QI��.��F ^7i,3�}�t�!��<-с�}[��J��S��#VM��K��2��a�ݑ#o�ހ
�'�����8��]s�ξ�76�gg���N�|��S��K�O ��o�=W�\魼H�U@���y��~y`���F]�L:l%�2V{�$K}��u���P��N�A���+-�����������i������֒�&v��tP	�@�p�M������ڣ��\v���w�<-�/G�$mO�|(u���>�ܟ��3�6�S����w7"���d��i(���/݋������kll,��ZԊ��U�S��p���T�4EU�?j�� J��ѦNv����֦��Y����WeO�i�k;����k�����(�jPI'>�v� i�gh/��w#z	��=x�,]àaH�V�]���_�������T!δ.GI��"���Lt�!�ۡ��y�9��PBKT�I�xZ�6�Ȋ�k�@���`�`���N��%�cl�����C�VrE�����Q�&9��ۼ�	v�Il���{%��q�nk%G�u�ʪu	����#Tc�\K]�h4&��_I~��/�W�ASAN��v('�����oe��~�
1뢭��e��A�H0�=�z���l.\^�� �t�%����@��� ���[2O֧��y�f���t=9�Ξ��h�RgD�1�i\�p��XȌB6�S�.)��x�tK������GԄ�sO=�/6�-��}�+K�"�ڇ��?p��k���̍ı�����?�̑2��~찑�\OUi����d|����c�S��U5�u�]0Wq��|r�,�7�~b�Lò�E�❮��港G4�TE�n���,���/4��~�Z��sӴ=�?S��V|�i�Y �?8C-($k7r��FFFVJH�\!��� �P"�Ÿ^���ר1�I��j��A'��Y�Q ����Ij��?C3���)m�F|�&q���sO%E�間���W�2���b�s��%5�UCS���1�*����}5�&����D�+�Fw(?�^"=���gտ��4F��5���ҽ�N�9��I��m�|II��2%�O�ٍ�;�޽-�Qi��Oΐ���OU��u�p����=����o�!ghH^kL�r��R�%IXp��<�����!�O�+�X�i��Z70`n��Y�66�&Z�	.B�Y�3����*h��0F������ϱ�7�|�[��6�n�4v�y��b�t����Dʡuy�2l�l�K�a�܇����`��>�G�z��k��3 *��-����wN�($�|L�y0�v|�]S����K��X|dH�a~s�j��kbX�Ӫ����C1abĸ�"�o9��_���V`W�:J,I�>�M�$���ơ,m���Lï4N$���z?L��\�X�gv������� �I�SG��H�|���(�쀪ТV9���X'�Ơ�����5挲��Au�Zr�ZR���yv�Y���[�T\v%�	��&�>�e"��ZQ����XY�(������fS��*n�.�"�Eh^*����(=MWptphҒ^���Z�y�7��^���X��CY�X��0��F�C�dp�j�@
��1�=�%�ɒ����gN9���W�c�cIL洛��	rJ���f���U��4��8|�gA�q";uR��M�}���M���{OU.��%�C����uu�q��=%��t�w	��*ӮZxf�|�V;w)5Mj�\m��s�q�d�~i��7�3��[ڊ�~u�����&�v U�E k��9b�@�}��h�����=*g�'e�=�6�4��@�����2�944�oab��Ig���I��i��z�2�b���L�SNkν{�c0����.e@s�5��$(rr�zL��h_LD���z�%�f(M�Eӝw/�c5	���ށ��ÁTW;P�;j,?��VM"o=ȭ��ق:�s�qTbELH���7y�32S��l�3eC��#J���TG�o��CC\����f��#X���m� ��%%��S{Ʊ��Ȧ�Ä�Ɇ$�����W������t�~�z��xW��%J���(�r�8��*h������ͽ�Dy�nN�t?u�q�T�&�Nk�"�P�����!�1377W��a��������}v]]]9f��H�0��G��VV��:M`����u����#4�8���)��3ќ!o�RY��m2��iP#�ac����N�u;��Y%��krVR�����9Tr��;�n�\#�vYd	�X�&�����d��-�H��p(�!�6	|�k��M�4��-���``���D�(۽�"A(�wi����ɳ��<�J=�����	���Y'S�lo��*������;��-]���Yo���Z2��M�+��Kk{FR�ъx�V�H�JN�ݻ��⭜����)�gD�|�@����"����Q�?�+��뷹\n��~����*�`d�`<����&�kG�\P��
�`#"<��yB���sqm�OE4����2�����2TY�r�Ni�B�w��o�J�?�5OFI<��s�˷�O��.���O�eT��"X�ho"��D�:��"�"f�e���L?�\�����䴨��'!qįh�|�?D[������yvc7Q��O)e��)�%�Kշ���g^�q�)A��%�$(3M���-����y�U/�yZZJJs	��XBcf���T$1Je�{d��ܘ���~6j�#(��]����������qq�°jBdI�6!�k�����qI��X�|�$�j����x���555�׎����R���=ȰV�Iy���N�_t���f�s�\���ڟ��l�7<��貖��Vԏ�	ԣw���c�6�F!W$�m����p��]�&�Wj�C���J�tel��DKօd@-q�����C���"����C���$l�b��r��[���L#X%��r9��U`�}�D����`t���(&��[ԥX2�z�CdA���	��W���)��{3�v[ٝoτ�ƃ���3D�ǜ��[����8"d��Qo_�ײ�ں���~�e_���p��8�p|����z=��[��o��}$f�pU�����Qm\��E�6`�ȠK��:�b�u�P�\��K�1G�\GnFĜ���_M(<}A*ݱ
����U��?������&օ.�By�Du����F���:o���֯�����cx�8�O� �[��P�l��C�z'�^�=QJF�D�넢 ��/���0�1�r*�S��S�����>�и������DF�-V�:F}eY�Xx�{�A���-�6:���j�j�p=��Cw�����(�5�<g�&��~�w��V��#ԟ,��n���$�K�Qȥ���{��z '%�+��zZh�d���m��h��n�Ih`��\mHp�#� ��5�O���K��ވ���,��{����r��E��	���
�!A]�H���FZ�<�o�Y�ΘQ[����y�|.��R_���t4!�Y��y��b}���ȑ7#�V��k.��[�"��r��#��%��)�kG���#bioo���^�.�:OM�7�J��DQ@�!�-j�s��%An�(1RjB��7�����$�mK�����eH�͡��lv��O��j�vF)_6˧���>TF��o�y�5�~����ˠN�;;v,���9"����[N������J�t��Ut�v��`|����N�.	�yė�B	i�'�R����̴��t���D�zW>�~�x�P(lՔZ���%!�]RF S��g�щ�ΐ�<	������H�����'��G1;]�!T���')(v��יh�*�tQ���&_��X�O{����過Y�֕2�?�;��r�djC7P5�5�(ʵ��q��?85O� �-Y��M���)�^���xH13�Ǖ�=��������؆�4nS��b8+g�o9�9�)fh#���%�[���_<��gЍ	)@�9g���)Ą� �õ��YE�갅_��Ox^ I(:
�"H�����=�ë�r퇴[��oJÏLf
�{^�^�r������<�!��Ƙ����j�JR��\1�%�~��gup7�A,b�I��K����s/V��#~�~�&p��E�#��;�i�Ԅ���#��~� �.�>��x�׽�@�y B�ie�I�����T��V��<��z9���A8�w�(6�{�ՄSOY��w%��v�=��ۼ�U�g�n��@[�?Zrܾ�"���`֩C-^+w�g�(��8�_?Frn��	�<v�tK��X:a$X=�k+&�"�����LN���Q0~Vk�/�21����5���w�ʵ+�	�7Cb�Df�Lie���'�!�Rpْ��cפ /L�5�Ί�6}��Q�u�%r���NN��萷�8¿>li9�������"�z�憦��z2��g�(kK�]�*��Y��>���H_��'�uے��#��{��S�jB��*,������c.��j��A���P�7�U��c34�_��j�Dp�u�C����@�\Ǵ���~�"THّ]�K�	G�{�����!*����)��ܽjj,�`oo�	 Zǽ��(ĨR-��»y���"�9��������i��n"�%8e�%��"%%%�qJ�o�_������P̢�~b)�9���"ەl��ty<�_i��va�[hÚ�r����~�U��������z6��y욡�˗�n�1��$� �ju� ���֒�\�.���<Ra#n�#Y#D(�I�_�N�Ԑ�N<��X�M��Rt* �ҕjVۡ�<�N���(�qC�k?K��rqee�5fG�Tr*۝��W���h ��tP�zt��x��)���32L/AA��a�[}��ک�P��@n�Q���X�8�s(y��:� ��B��goQ�đ̪d�N+�	��X����l���x�]�܏��5���@F���')>�=�����y���5�"@0�r�A� X@��i:�]�3������(��0��$�!�A�����J�3���[��~�)(&�&�6
'I�r9��<�evM��Q�����e�/_>���K����.�m��ur�U�K�S�����9�__�?\�5!�,�]�r�X�g6P���Vm�߈S�xo-��t�Vvיڍ��^�����D��jFzZ5���j8�uM
���䜈��@�1
ـQ��2��]:S�I�ѱ��ԓf��j��o"*d�\ ~r��q����j�:�s[1iH�x
>�+Q�/��ȿ��G�{(IM� �*�B6\ܻ9������V�vLN�7�������-��M�=~6�}ͳۄ�E��@����.k�*oB	�Y�,,��>�/�	�쯾3A�h� A���Dm�E'�b/g�Sܙ&=$��z�Y�,�>.j�Fn=��Ҥ\e��"�W�kį$�1��:�����)X��"tN� F��f���ꖢ ��:O��>���Z���X�r����/��^s��]��P��\�#��=�{8�i��{�$�~<�λ��7~��<d��۫O�&����e�O�G�{Q��=�u��v���U�{-��7���3��U(�9N9�v����1�"ף��	*�w��|�w�������0k�..�Y끅�!��n%��n, J"%5UKNN�ƽ4��(3'߽�ʸ����u?�u���~H�/X>���	v��N�ՒPns�'�x�;�@�AM�)�ދ 1&S��(-���,�Ă��A��k?���,��i��hg�RL�SV&�_���r��h��"v����F�y���(��i���:���rDkk`�wtoH�8����Ī���&����l�n&��~h���XD����PUy�	������ce�g��:���I��K�@�(����%�a,E̺�G-������ߠ���g��Lf���F9-Slv����yE����A��3����'�̲9Q�����Ch�_e&qZ��V�z�5��/1�����%Z�����ה�.ҍ;��>��Ri��Ҍ?ˮ1���a����>��z�@�I��T�S�+��zk�v�<yc%��3�������Q}_�mv�Rd�w�[t����5Ǩ��(��J ia�Ĭ�2�J-^�:~Q& N��i����8ik�_�֙u'�.�����5a��w��V�1�aw!{�5Hk�]1s���	�S执��?~����g4�`�L�offf�	�C�q�\�bC	�]K]n&�R\����گ�6�&IJiyw~�oyĪHCZ�M�q���:`��w�O��R<w�U�ps����V�9�������b��ݓ�ĠW�������í7.c/!$g��g�C�4���g��w�m�Lz�5W;w�;9̺D>N*$��׫u����j�X:mz,j��ɗ�a�g���Z�_v��IN�v֦\� ��_�����;��v@ʿϮ��O�d$�NNo�ѯ�B�:�s��ū�.�r�ϻGK�&�f��=(6vin{�C���f��ࣜ��M���{�7��g����������i[_�Z6(����!�5�"�E�@D�@�~�}ĉ#��3XQ@�(q4,Q�FQ��o̍>�R�7��{��{���~,���2�Ӕ����w5�j�
}��D��=�!��H��eR�R==�H�Q�/ef�?���nD����|��_Q���<��!���O����u�Ɖ"��~��:v��Α(v�U���&=��j��,\qL��)�4-qJ���`q�:z�␈��� E�
�Q	a[�l;����*\���A2�ˎ�X��N(���u6m���8��bVֈ;xZw���׏����^���θd���p7,s+�5��'%��8�U%b�8�fr33��!+�Q���[&���1���!D��K����#Ʌ�\�o��a+@[�˵�e�da�.Y	���X�ҟ�`ہ'oWh�-T���*ZNNNk��J��9����,\�Dת�(�>U�Y/r��p��4MF�=�?�|-vlԏ�U��J��!'w�J�w�Ĕc+�%��/)»8ΐ{�J  ^ 
�>F��_l;���O��:@�BZU��w��ۋ�Jm*���Օ6Μ<�t-��LƭǞɻ6�YB����X�
�c5�	>�K)�Tff��8��:��4��z���٣��@�o�lNff�K���k�\|�~���Ɓ�V4{R�MI�߸q��''����0���au�K���@�%*f��C���$��������t1�({����3����>����?�Fg#d	9��F_M2������5{y�o� o^� �ݭ{Fă�'df����V��H��Zs�\���ɠs�XK᛿x�~�w�]�C"�N]�G��-��eӣc�7�r�Y�jH�,�^�?�N�͜����!�`M��~��u����~�����Č�Bg5�3_���݇����W �����๳|w<�qi?���Gw��n&���?K�ea��ZW�L��f�k �O���+�Kܔ���sY��wtc��#�1O R�@�[G0�o��A?(��V�g���.I]t�#���[��E���L��v�&��1pk�k�z��	4��Ix�����O��V//�ALL9�
W��q�;_��U^�+M�������l������[���7�KJ�&��+|ޏ�� ���>��AV��ݹ���CD��_��v����"{ֽ�i��j�b�.z��E,��,?��
J�/���.�u�yw�\�?X��!nT�2���{�8ՃD�������D-ӐW����n��AF*�i)��lȝ�ַ�9����<<�$V:�v�JP�x�-��y���?Rec����u�_�RH�dK.Z����7�!I�H�v�����[����l[�N���]�����>���t���\�="׳�J�mҷ�޽یΠq��v�ƃ�6��c�ݤI{���Y���+�H_�u��g7��3)-���mA�J[Jcq��$Դ�k�g�����}Tԍ��Is�Q�E�^��F�e�>?בF==g9��Az2��p;�m	K�Ŗ��糥�7 �lG!���?�2��3<��`���t~����D9������l���|+��X��+�O��)`M<d��<^,�i][��	�RZ �FOP�̟|||�YWH���n�D�5JT��[!Wc��s�&v�%���gpLS__�J�]
������NG�$� �A�S�b�����u����nz�+j����Z��!�~Q(�|-�`�f�6�7�����~xH-�[Q䠦��چ]q��85[$*�I*@<d7��9#����(1����v�$0��DY��[�f6�p�b!��1��� G�M?/{�RÌ�I�Q�)���H��2���N:R���|��e�&q��n���?y�~}Bqa�Ǐn����z^~8G7B���.h��R�uFo;���f0�;"%�}H��:���E�*�����,f$F��U��7��
�u��@����%�N��O�+:21o2M;��7E�����n��n�g�u��r����v����y8��k���4������C��ʬ�&:�[�"��� y:��>� {�b"��n�]nۑ?3.$O�L�~Ȕ�O��xU^Y�c�G9��ƭ$��6���[�-�7���p��9x �U���
�������]���� "�&w�o�<$�`ڜ�����y�Ђh������
��Syi�K
&R'���Č��G+��L�m&c�-+�|�6���̧�F.=���1`���JP��¦�>I�V�av����&�����o	�U�ڎ�R��_�~��<=�@E4&C��i��p��a�j�u�y/����|>��v����iW� �𫦙�d]]4g1�k�Q�ێ���x���4���t,�~�Dq�F�t#�g���%5l�F�-��ִɊ��;T
�����Eާv^��7�x�+4r�P˔��h݅ǑCX�Dt�i$ܘ�Y�����;��j���;�<���J��1ߙ�25�7��hX�����Q�ω,�c��5��|>���G�:��{Ď�Es!�cSe�O�(�d<�]q��{䄋����.���%K�78>n7�61��qW������u���B��3 :��Ш!o�k^�ΦBfے��q�.d�3�M�M�!���ˤ!��I�L�ސ�~XM[�m2W�2�ʳ�	�O�>�F���I��b#`�
H�W����i�*�ã`��8��3].���M�9���MͰ���
��^��a���{x���.:E�;��%�P3�\l���0�I��m�1z��v��jժA�kw�r>C`p�'Y��d�|I<�������D�L��
�ƀ`0�Fz�Zm�I�+v�)����F�O`��YO�2����t5F>j�F=�P�2���(|��?Ě���6\ugG�ye�i���ш��=��"$�a6����� ��5���oY����#`�|޻p�,�oH�0J�VyG�C��sS{<x��(|�P�]:�;��b[[}6o~v%a��IW�q����O���������酹i!M�bz��L�������۰�g8m���]����
�5z�B��%��H�0����A6B���A �Y��k��r�,^=����Si��◔��q�#c1_joAmU3�'������33[V�ܾc$����)���lm�S��[�m�2g1�Qc'Ǽ��44���D���uq[R�c����Sxu�X��b�e���m@u,�m�����t�a�:�DY2�'p}��Qt.�`��J�l$5����� �;<ǅ���L�&<E�p���).���]1����FF��l��E�Y��v�4���f{���GqNGtR'·Z�`yH�-�s?r�X5�h+o*�	
���5xֺ����&���&3i��?Rv���/�����f*J�Tr$�p�E<$���au�v�t�^D�9�3�q�� �e��[�ϔ[uE~�<��(%����3&f�2�}�mSp�v��w�ܙ���9�ʁ�~E<���kܓe"���^$������^[Ϧ"g+9!�_�Z���e�12��`���z��`����6��Tf��0��A�`��P�1S����mY�z�]�$ FNsS��UHa���f�X�:���j����r4���utԫ1s`_���n5l+X|�j/q��߄���2uȣL�͚�F��0����l������q�]�a�b���&P�'~��E[�wq��	�T`��uUl���ׯ��%���R�D@�ϵ��ۖ�Ӏ�1�7&������F�m�
xS��� 8��V���y�zL$��S�0<��I�Fb�33��Uj��1Te4�(�vj�"���+3��c?�J6��W��Axq��H�Wf��Ԅ��]�.ŝ[��_�-��= ���\M%�kyE�Ak�K�������.���������&��:؝�?Lh)i�;U.�}��Y�����'�n�[�D�rO¤��6���.q��vu2.�-(��H��(��=�g�ʹ@��l���� ��L�tt�6f�'�,�~�p}5b��JJ�����tTB�[=g����Ss���Xﺉ�F�b1�`-	�uu�3���2�Z���|6b��� �=��b^�*&�N��B��<�ሒ7#˵���?�%V��ӳ<��T>l�Z|� Hј�e���kF��(em��8v5/�k͎����(y6
�3#v��D
��^͎�#j�yYYY��P�䐑R��s��
S�Ջ�U�7��[М#YmhO��gΌ�c��e� ���:�NDyY��˦MÅ�ù�\\���m��- 7mA�H�4����Yr�y���K������s
D-f��K��6	C1(5��׮�KblFn�n01�|��(%9je�6�������^%!5����X���D�+�����,ᾤ?���`>K�0�m,�s]T�K8'f��\�tZ�H���Bz�%��[�ʶA�n�c"r�< ��D�%6B��`��S��؂5��E����n�^��~�SQ�5(����ŦBC�?#��s��G�����Tnʗ�J���pu����#[�(4��Ex�]��j�D8�>³�lL�+���"�h�D����|�B�������D�X��P�������9a���n|We�F�da��+��AXm������@��_J���=1��]�[?�g��^���� �}�����.�5��=��y�n���"5ݲ/S!��}��m��kD ��}���DL�D���CeuU���kK���;����19ݥ8�@�-�˒�,�aFM�lCi�s^J��Ơ�{xk������O��<�������~4���.�DY(`s���s�Cm;1ziE{��en  v�-WZ�TZcrB�1-��`\9'��hJ������OR<�ƚ9窐����*Y�pb�E�^�z{�J�궉�u�B�9�,�_��\�}^�q�m#eo�$z�>	6PԷN�@ّ�괤��H��j�:�e�J�$X�)h�E0�8ÒF��u��Q��qZKs�xQ壝��5�WC(/OO�4F66��?{�v���N�nlf�a���1�p�4�X��ȇx����$��ppuՌ�z��H0bl�>�Q�),J���ˏ���'�Ho5Y��Bf���`[���z�mG:��D|�َRݏ0��c� �P�>�*�CL�
㊅�$]^a���t�����()��i?�iN�-��c����?~r�.E�K��� `� �$�ϟE��vA!r�2�l������j��e���^�N�M�kE��ҕ��T�YIW78�'��s]����?�-�;mؐ���E�8O[��>�b��7!�o�ݾV��յps4�cmŞ��H�ZQ5��� |!��[�;
��![�c��6PU~�8��u
�U��S��3�Wc�����x9ZZa���k��������e�����8�ۈ9�o��9��h�Y؇��uA��ӯ\�rvس�Ѹ;㳒�Z������~��ne�"f���þa/�œ�*Fg���N�e��:���;G+�����vV��ʟ~�G&8�=���z+Ȟjh�
�m`P�&ƫ��ܧZ\�{B����X�H���s��I��A2��qS�_�ό>Y�'@;S�ѝ�Gh<0�����T�8a�'ħ^�6J,�c�wx���v��n_'h���K�(�O}���aQ����;��ow@��B�D�b�q�+��P�G�޽����E��UbZ������4�z�  �^ 73�3�#�ع�7|x����F�i�`�zM3ng�eБQ�w9�CbdZ�q����~���~I��PΓ��m1��u9g�5���	��R�B�<ؑ�����H�h7��u�w~E�<�� !���$Ƌ����4���l!��jo��GSccT,{x���)O�PV�$����q��}�p�o��nᎧ�!Ğuqv����Z�����s������+�g��f��ƺ�k3w�R�� .5F�������{�"��nK��d�C���5��ëن��Twf�AᑶQ���X�Wz�Z��w�T��`*o������!�#�p`�q@��7B|����ŋ����X��6��T�Ǉ�ʅ�==�/��I�����	R]d5�~�s�S��*G�,մt��Ml,���]��Rn�i���x޻� �@��(xO�$��xC��?�
��+N>����d�F����lݹ�i,fz5�\���_���DBD�f�]����L��|)''�	�JyS	���C�B�
��|a���O&�4�a$�}��^�IQ'����J��͑�b`��GR�>�
wU����wt��p�X���4v��e5Ht��*?II��7�̶?Pz]���ll"�
h
�1oY lTg�"���95ƹ�<`�@�^;kv��^W�M\��A�3n2z�Q$�?�O�*Z�SF��7��4�֕�Sl�8���_�mt�MCv�~��{m��G4?�}�e�O��opPݤ�C�O�e顇��#�Wv��?��昋��	�_�1QD祪��?���dD�fj��t�~8����|��n��q�>���u��ٔ
L!���AGky�QY�ME�e �����砞�k}��0W{�-��XJ>�n:�<�=�p���O�QB � P��d�\��q ��F�J#[�E��P�y���%ާldz1B�.v,�_T鈎�^ɫ�������ZЋd/!�-%D�����T���;+w��&�Ֆ5�D���έ��Q���0��>�v�Þ楩$ܔ0۞�"N�֜(1E �1�ˇ}}}�A>����0T�,�!�@�v�?6��.�N��%*$�2�
���{�2�@V�;�&|�tP�h5�/k�����Բ,�D��N�z3&��������Y�������B���]$�Ի8�@8�\Z�6Q�>.��ZʴH9����Z醡�� 3z����Ӳ�aT�n��ea�..�,���=d�x�߇�_6�#��y�N�����%�5�`4�����1�j��K�=��;7�B6>^�7U����y]q�8��܆�BP��ۻC��3�!�_-@}2�$�ڥ3���&�ɖwJ5WV����7�c=��K}F�j���o�}[�D�w��7� [�r�n��/B���F���d��f���p8�����= 3�σ�o@�	d�#��Y�%�3���7\��O���u�Oָ���^mn�h���YVh/�_�
T122��ɷ��A�f��{�ғ~��m?Y�����Z��+�I,�U=K$��ϴ@c7h�B6}2�&�q;���>��w�קԓ�XZA�f�ɪ��U�ވ�#�"y%8���ぎ���l;���켼<�j��&1�`�2�oh˫��^�k\�Gf	��0h���#o��vY�u�l��3h����U�����V-`��<�_�~��e/�n7g�[�A�\��í�?�]����Y�A���i�?(q����a�d���֭�Gy�4��ڞW%�"�;D��]!�;�Ʈ؎s[E�s���婜e�Rͱe��QdJ<�����ib�f�L6��P"@����b�a���]�3'OP�� ��G�h�c�t���Q�����q&$�R��`ڌ^;�^���&ʕ�@���S<��u!��?���|5��<���5p)�?K&IT���Av�$����o�H�4%�f<�S�[��9ΚU���@����7{�K�^�Q���}��LZ���^���r$��|v�����i�j���4�s��s~��4<�[��^�7��L�>o�(CUC���9:������0\/%;��Ejj� ���0X����>>>swf�!����կxx/�3�;���P2�zHi��Z^�܌f������˗��ə�A�gO�xդ�m�~L�� gr�4�t;x\K[֠X�s�2 �:900���; 37��v�$�9���S�6�վh��+����� ���ՠ7�������2u�-�ϴ�8��a������\�ja���0�_ET��s�%Kzy���<r����R�UM�{�Ǧ�9U\�Z���D(=��q��w��/��I��!y��#�)������Wo���Uq���٢_9��?PK   ۍ�X��L˪ x� /   images/68064abf-29c0-456b-9754-5c6c0ecaa6a0.png���W���?��6�(JH���t(8�A��J�0" %ݨ� �����2t��:�0"1"����kY]��������=p_���G\�����¡�P(�!ū�7Q��%(5۾=��?N��?������>�L����^�أP,o��)j�5��28��8���qp�u�rvv�7���7�e�巹o=%ɈB�B)�^�p���s����$�I�U#L�?��}�;�-ݝ7�䪰�}�ư
�m��J���N�?Kw�W�7�r:�e���"�S{��w/�)�\�aO/�q7�=z�/L�����W�.�����'i3�v���,%��M�h�X�d��~��A�������������$w����y�,�B�mT��m{�Oճ]�aT�6�)��#4�#[�x^�ӊa����,��4y�j���4�~/�	�c4�4m�~�a1��e٘�~"��4�z��x��	�J����O�y����3+�M(���q�<�(�d+�T�s��O3G�Ӝ��?��N5�ڸᛲM���4D�1�~ǰ��`�gX�Z�7SY&=����Rޠ^?d`�5��~tt��&�K1,?�f`e����s��wG�N2u0�a��}02�L�!n���Hk��w�~���Sd;�˳{�P���s2�����)���s�/�5�є?�0�����z����auXC[���֢�O�ֲ�N���=c���Z�v�NmCcc.7a.UT����ZT�X����콬���hᰫ�7h��sy���*a�B���}�(tx�z):�BCCy�q�Z�Ŝ���pX8�m��NlF\Z@�^�\�d�6�o�f/5���#J����G󮃃�Z��U�,`��=�(�Y@�ԗ�F�5N�9v�>�̹s��c�(!H	O��ϟ�s(����~�|N����[��ɮ���3�*q#Fg��{���G�֧�5���Z� ���V�����e��i�O�@˱��r�g'�$�Kx	��՚��^#���1������Ԉ|�a�����v�͸�u���;t��7l>�7nߠ��e<���\���xS��:w֗&3Ţ�{��[�*��nK6�̲�;�W=������$[e�Ν[��x�������W�+�y��pXg,�IOvA���2y	Cr7$��֛��>���Tw<���#������Ԫ�T�Φ'��TvM1���O��a!m��q���y5e)}x63��D�0|bRɇ���:u��d��~nKH�%p�c[� �����W��%��Fi�B���=<6�~+�*��|��l���+]N�5�1��@�g���S2�Q:�);��d�Y*YV�5������+����F��RfX�2�w���Ywo����N_H��A�Dv�R�a�+s�.��Z���K�O_BYᓙ[U�ll�u��,�ʬ�d[�%w��0��`6/��
[��<���.�������^`PP_x*Y�E!��_���Nt5��0�P����i5H���aT4�ߏ	��]o�%�G��33�v�q�x7���K��m\_��1r<�"j�u�s�����<_��BdU".,q(�C�v����%D¼��W+!��9p��[_��$ܗ&J3��nhdk�����v�r����숎�9�?����ڢ�Gyq2.������G���$��w�Њ������O\�nGg��J�z��|rҺ$��nE�an��b�ϸP�O�[��JĶL[��-�.�����N��Q:�������}c��#��%�����'�I����ù����:����\^��NQ�	x�u�B]�0���*�*īax��!�\�7z�F:,
�\���F,h�Q�)T�����0R��M�_���D��:뀎�[��f]\=9��f�)n������O�ͮ[���W72;s�����
_,���\�^�ȕ��H���z=�g[{褻�[�QfG��p���JJJt��N�=^��ř�;3��!�'�,�I�����
Im+�]�n��tِ�-մ�\..���1z����K��̆��k볤��U�cqw�͹u��D������'�I��X����y����6"�dcK������ݬ���l㶁�7hܙ> ��d�x	^h�:����)��`����I&q������:�s��ӳ���}�zS6[+mU�C��m(3��f���̫�GYsP�v�Vt~�e�����}���0�������5��v�9Ơ��� XV��=#_+9��w׭�l��b8�*�ފӞ��b��~=Ơ�;��%���S�����?���x,�����T���PF:�����6�faK�i��m�ߺ5��tAX�u[���K��4ߢ�&��{Ǹ�g(� Uwk��HK켩ӿM~�ҰZЅ���***YV�L3�S��H�����Q����yyy���5���Z�ҝ|���y������!N��Gw��T�h��;)f���zzz?����|�]]���L�/5sTf�^c)$́�Ћ]\�s<4�S:f�KP<�gtlƳ�Uu|�d\H%vCe'+"�z`P&'&&rY%��危�,��a~��������Vn�7��2��S93�PZZ�"6v���J����gd�OHH@�(j�ښ"@��o�ڹ�رcR(�nS��"]+��%/��ͦ沃�Z!V{{{!11��;�c;+��1�j���HEM�������f�'G �R=uuuo&,������ܸ\i��K#��V\�3	����D��x&C�_hW����y0�x�%��\^u����ʽ�z�kt���E)����K���þq(���p�:::~�j�(4Y���Q�10�=��3]��=����>���ʒ]��88
W
f�Pw�(��Ͳ�/��۷��ZZ
t����>%%e�������P�{�BU 0�<���o�2�)t,{sJ��27����-�BI����#-���f&w��2�ԡ����ۇ���RU�o�on�+��Rj
�4�f���`�u����Y����f�{�Y@���?F�1���o#;d���^�i��2O|}�>=�Ho�.��l��7v§������&�An׶fTjy��kJT�)��iiI��;�D�}��������;�?��H�Fz�ho�����Wj}a�>�ը�j�	���G'�$`���H��4Ae�C}�x����F������8l�̏:����۷��;�.nq������)�@b�_��nkz�^�yM��Ϋ�K3C���a������%8[�X��Ʀむ��FPD2Q11.|�̠3������f@���֮ xe5�F21-�H���G�C'op|B��LH�Dp�ί�In?yU�Y��:�GF��@�lF���8������I�LS���i���`����	;Ϫ�htz:=��u�^;�$>M��G��П����u� :�KQXñ���nm�\�rG4�hZ������EU2[J��,��,V������:�����y�W�.��Ed�S�4�����;������׍�,��9�9�Xxir���ӧ�3LPZl��_S�664x���� ��<�+�H����^GW7�����\��Nu�f�\hx�̎�rh��t�Pa��VVV2A�Ղ�j �)�>���� s2�;ґu��z��AH���� ��%%+Ւ[+C󚍨,Z(�s���-n�:۽�-�c��`�Z\ �e��Ί>@�|.s���S��t\��?�L���efI��k
��0�6"����9��*
0,BXL��P��c����9�����y�/�NNf�Gʹ�L.U�v��H		�]w���(544l݂;�F3��?�2���<=ƥ*�ߝ�3:O�<����h��!�,a�iJJ�2����j;]׏S:�bc��\��s��V�p�蛻<'���3���s�0B]�=ō����m
uY����~(�Ǳ����5�k��Z��1����[�p2����x裙��+�4�&Z�&=���U(l<��B[z�
��D�	o-����D\�^�3մc������>���u]$�݄_B���{��C���0��WP8�LY�&&&�]�2*a��|�"�.]=m���g?�ؕ��U6�E����"���&��i\MD�� �ʱ#<�lq�K��v�ݒ��zZs��x�~�C���V+d��ʞ���� !��}~=Pk�o�H��2 ��2��9��j��r��TdϞ=��Z����B$��A�B�yy���V,�ɓ\��w$ !b�R7;�hbn����}l����ϥ�fKKZ�s*��7���C�ƾ*������o�@�����bЉ��g�ĉHH���	���q<�o�^� 7�p#�����g����-,�r��K����df�� EͫB�QT�f�\?1q����0Q�v�؈���v>�>�Yq�$���{[@^�HU�b���������(�@���A�������/H�{6�رE7}���yX�jX�P-�_>Hs)@	38�K�V�tV�9���?j8L:�v��'#�*���wd��!Zՠܩ�G���ܠ��l������t�V��]��Q_9�W�=~�7N�(��x/4��P��.�""�s��3@�F�Q�������[���%cG|"�v�I�/�w���Ƿ�2疥t�khKR0�������9JDQ��	��<�ds]G�n�dg8�txtz� ,�Ԉ�K�bؽl<��� ?ೄwW�x{o?!������j�k�wD�����������`���g�:��ި��aL��X�T��:��e�����j�ų?�NFZ�9`���*�����G�-/7&VWo�m���8$�;Aoʃ��f߉���K@T;��6ĿG����'�=$�K�ָ���n�4�Xh޳�̩��0J&�$��O���`H�={��dL�5 �\�ϭ�@��g%��%7� X��{2u���(/��cD`�q���#�v���+W��;��{�n���ohjR��`���($%ŌL�اtq�1����p���HURE6$ś}���{�i)ۯ5�'(li`x��� ����c1Nf���# �Vf�@�h2dK�4�� @W2��Y�53c����L`�b��ц������F!����BL����B��:�+� J����.�%
�(�(�	���,��쐚��s��h��`���i��+G�?�}y�dc� &=c~gw�?�n���2I8�3K�Pa�wZ����=�e��Wf��:��E��F�xqW�Ō}I�YaS�*���^}�U�B�LjƘ=&ON�䔰9M�3w�O>�Nj{�޹�4����>��V���ƁZߡL�M���f��a�)����p�6�D"�#�H���RF�[ì���tWԋ��,�pkSSQM�y�H�W/�]4(V�ِ>��2d�ء�~v�k8m�&�]&��Y~l|LM�VZ~�՗n�_u���
�Z6ߙ�{���Wvʇ�#�$K.������yI$�4�x�)�ƫ�4.�����J����6��9��kkk-;NG�r:83P;��$�T���7�~�:8l�eWҵ��@E}��B���](C(�1b&A�{�dvl�_633JO���x9~4/��ki��������ji0���L�3�l੏�H��>�Z��l<�����Svf��]�5�6Dێ髄����''�?��ZNu[�[,����$oX�YX�(�S�6F��u��o��%M���1`���'��Ѕ{�,!h����P��ϻ�wot�X=�	��1��E��\Ap:�ż˓��������Fi�#�˱�>�O�������\;Hm�`�ET��/����ӧ?��kr�
:t�^S�@���,A5m���V��[>6��<M��A��"�a��1��~@w�����@ot�K�'�K���Yߙ�>l�۷�`��g�$s�O��ved� |����r �/㵽�����A�=�G.G��ݧU¾�+ܷ6V!��p�aI%�dsFΠ�����Ƴ������?��>�c�z�c�`�Ad��Q+�6d�08��>��m%�&����Z	X��q��:p�nN4��H�$��?<o�8o�NT�l�v�Y��/]��e�̻������qs�_k�̼�;D0��｝�KJJʮ�\�,��QT|�7��,bQ�"������\Q\\\�b{��t��{�x�	�u)�'�25��y"VgU�W4ac�SG�>`�a��ggj+���O�b�K��|�oŉ�y�?�	x�W�1���W�p����J����������a�]͑��.c�i���l���{��G�S��P��˰;vl���pݷo�ϱǣ�7A'��,s��UVŘU�(�B�KȲ�3u=���mY�1�0�bce�A�R�����T@rKL�ILW�����Y-�`K�\�u&y"�)�~�D�._N��(z&&�"��42����9���5�@B�[j����G4y�C�e��aV�JpX��GZ~��cS-e]>Y�����3A83��tUG�{���9�@ �|o+U/�� dW?ᒱ���AA��U�tR�����}{�n��B�쁉/�<SU�S%�K=&��/*W?8Џ�؞z��
�k~7�2��<cP��XI�?�_@1>F��Rfojhl��!ږ�ͭ��"�i7X��:~���d"�����4�w��͋s�X��^�9���K
q�X�*HS15UUU^$"|�_X���ZO5�5f���X�i�	��+;�D�B����S��(9���|}�wP$~U�Iƫb,���!zz��aQ�Z����f��Wj����F"Wy�A� ��:ɕ-}��s�z�U�����t�3x0Ϟ=�%�y�^y	�:�SJ��2��27�083�����ԭ�����FE�oA	�"^�1��YyX�^��鄒�8�A��_t2�Y��������i:�u(��n�c�����Fײ�E=��\�)��Ѧ�M @���+�;�I��#�p�K������z=��f;��Ν����i��66<zݧ+��}h��̓[!��4����Ѥ��F��75�ewMM�����{��mXfwX�9��I��Aq�+��f7Iۛ?$ݿ{�;�3�^1��b�Th��O�;u��իaS�r��A��*�D���i�'h�ˏ\���z�	u�o��2I{��cU�Zg�x��W���4��W��L�وW�� �@5��gv�m���o޼)�
�5����4M#��߿?��ò�s7���C0���)���q�3�����O"�{��fs�+y���6�O��%�Q����NA�hck.ڬt��J)wK�%�k:��[�Og��w�(��6��Y�0�^C�I�M�VG��
�'L�|����"FK�}e6\�G�e�`����9o��yR]��l�a���s�Q��)�K�B�� β�%�e�t�k|�&͐��߇~�d�:���.�n�kzY>�i���N8�O��,�9y��#�ɐ�
���S}ȅ$�07����.�-[)�H���;�2U���+k�(��p����rǇӷ�:x����*�����ft��֧CB<'Lق�E�/�u��r\��r�y��a>h�ٕ��V��}���<�(�0�bX�u����lݱ6�C��C:�5���|�������{�7���}�{Y\NI��� ����P�0�]��\������>}����{ Qq��š�UeC@nu߅��u(V��eQ��Qsx�bŸ������/��͖�gG��Ff��<ς��:����熸U�BQ��|Y��Δ9��cmq�������(�2qa̺�e��lh�-�om��ovvve�u{�s���O��z�����Kz�i�r�{ҙ�����e��eYP�]� m$�o�
�]��5Q��i>
�ޕo�r�8�{�#�0�o��fX&e��{�kHj�U<������ǃh�ٲ�J~� ��C�R5n��{S$�JC>�-��y�T�䭉�֭�&T'���o�@��tVsSӆ��<4�eP�^5��r/:G��n��e������m����y��_��$������q 4����>���f���\�ґ���L"ƛb���=�$[�,��u��8�M1'l܈у#^S#���+CS��Q�#W �eO�{�%B�˳Q�&W67�+�>����d��{��:���5��jC��N.%���8��K�7�?��ϔ��۹�#1�<Ie�*�v)����7k>��`CV���Pj��GGl���;��G��!/PG�.	|�x��h��"���J�h��}հ���N��H���xtQ�}թ|I֮a��鞑aM���
�e.F��M�s�Ι���36ټ����YU��ym�|�+++�ޫy%2K8�a��nQ<CLS�677�h����������K]�������1SFf����RMڭ��U���V:rҬ����GA۴�QI�uԋ��
��@$����D��)�ɲ�f���lW>���ʁ	�Q�F]�5�a�O����Q�yӋ����,$0�Uz�bRRR�4�w=�������7.��Q��lu���jL�z5�kk>�0�!��޽���@V��(�fFf��Q�%J��m��S	����;�+7/%��02�TW�����#n"H2Ls�����[���h"�
)�TU�#%fw�'x����LiYYٲ��[�]�-4������!��:8MFr>�TTT-�vOѭ�ځ��]F�z6��rrr����J���SQ�b�s�˗AN~oo�7����Ĥ���Ugs�������]N�����{�,���m�����ZM�β��a�\�r��,��r�U� �|���}^듺��ql���	^B{��|�צ[i�u��k���^ ������yv�Gö❴'N�I�����P���Js�а?���q1T���ڨ1�Y]�)Z3������J��+ Ao-U�`2��S?#%e0ޙMk�2sk�C��hg��a�+�xe
W;��e�LZ}{��6%�Qp�]�-��9Lb�䯝l�VWOҳ.�RJU������_q�{��)�1��.0~��Bl�_�Ij_�]j���ܞ�R~����:E���Hqqs��,--e��%r@b$�|�ʅ�D��lp�)N�}�r�Sͬ%F(�hW;�Xh;���p���Z膷kkko�LM�+�E��y�i���n���G"lD�����	ޏ�ν	��~_�cS�H!*q���9�~P�ԑ�P����=E�N9XL}�	''�-�۾����J(�SSSO��ރް�h�7)���D�S���9p����-�/�
B�ҥ���Л*\�)w��U��|�v*7
�����������^=�[k'��:1=���t�v��u}��C'Ϗ"�eT@�?���b�	ᯘ�\�ة76>.K�x���݉S�.�*4��o�0��jjj9����5mmyF,��)w��|�9����Y�s�z߁=����(�ԥ\<u*�+��ÇW�K{�}�*���8��Iz�8�$8���.�WRTt�t�Zr�����`f���gh������]񣲞��U �^w9\���������le�����ј^t�gm�$7qe��do�V�΍	[q��27��*��$�}\6�"Q�@�?��Z ����۞���0W�r<�8NK��f���b�1�#T�=�$�G.��0�o���\�/��V�y���P/�%�|�u�o���V�������N$^@�����?���ڳw/;��uϒ�����u��EY�?����*���ɩj%;xI�9t�p& �c��
�+� �e`�ؗ��'�>�b�x������9a��h���`����Шe< �����:::�RR�I��-8{�l����j����iI
!g���z���̔#_�[Cp܄nT�/�Ua�TS!ǔ��A+**�2��V�so߾���gw<���G"�=�S�NrJ�f?>��jݾ?���nHK�c���&�z`�lл����kjj]k�����?���ʡ:t�謘���y��jf6��v��ϋ�'TSKk)�9*�{d�(��
�ӗa@���B���k�cT�~PŦ"+Mmm˵2�����7/��%B��gz��ޏ�����9{�xwGG� ��]~�v�����}tl�&�����f�m�:;E..��w��_Ȭ�)[���^j��_����,��/}�:]WN�{ة��G@uЇ�%%��lfՅ���Ӻ���4p�K����[��T&�	��zz�h		��� ���(C��;�YJה�X�GG��^D��R8s�Ώ����J�`�nq���Owk����-W(�~�f[:������|��ap�=�?vYܻ'{Llm}=�d�b<ӹp���#N��}�p�1��VhF�P����g\3l5x^ϕZ�N�����~����j�	�f}iR]��|,��ہ� �L�/��<�::%�C�LAY|�ka��X�0�>�U����hacIk�O��߮ ���[�����uQb�&٠��?�����2���ucr�6�2��n�|q��SiT�#�Z���?Z���?ߝ_a������	���X��£�#��?[;o�E��ӧ��*Oh��c��s{��Ѹ~����D� ��hT�C��YP���SD��t
X���db��PCP��s��?ۼ(�����+Vm�ec�K�y1��><�
��!�C����=�'��T獏�Q]G�E+մ���q���ж�����r'�9�S7o�J�m����)���jEh(��M'������L��gϮE6�w��$�5��B��a


��W�c+�e�<��BQ8�j�#���T�!%C$��3�B�WL,��+%%�5My�Ӑk���X��c4�v���[�U)BO�����>���?���
	�z��������N����0���<Zgxx�`>�*H3��f#�k��ILL�3�q��v}]�ћ��-}��i.���I-333���0���&3餓6`c#[�c|��@"����Hgh��Dd���r�=Lgww�v�HdNE=A���`&�z�b:��'[b.$]�r2��ia��{����in�(���߽��xA������Ōׯm�t�e0---��{j��
�N�n2�ꉓ��"//��{f���҅OE��,�ߚ��r�֗Bˈ�jh. iQa�DP?����l�#٪�����:�x�^^�^��>_^A�=<\�A��= ��՝^[C#K��w�4��־{�w�GKK�3�%�j=vH�dQ���� A�3(�-_�Ӗ^%�6e�)��?�*����x�_���"4>>W3Sف��A(�2��""�8��^µЂ�����PJ�ph��׀��V�-��Ǟ˱u<׀'Gb�-���ɧ����nsԹ/�f!@���Y � mޓcV���"����{�����R�`n�SC[�4怶�jb���D�K������A'�9O���]G�a��;͌�}��0���o�3��5o��%D�\(�2
��X������3HE9�������[�οH��ht���wTI�|���f��@�H���	���3�ȣf	q@gq��nd�[F�����L�=O$�]��r�ת��U&C{ 4�t�@F�VC ×�g�*ѿ堼�nTg�A&�����Ȗ������KA3�Pd%����;>�,/x��s���%Z��������վɕ��i_O�|���I1k;���QK�.-���{s�^�b�(Ϊ�����II���ϣڀP�\]]u���>��S�j�t�z���07--�]b��Yn��gĎ��S���%ai��'���uڵ�����&�O��N/���Mѱ��9u��7
xz���d$%d�f�V���m �<�o� {����c����և���Z�^xc|��������ێ��������W �8�ê��ڞ�E���W��0��ρR����D�E�َ�NS�:զ�U���ӱ/60��i�t��`�o���[���ɴmZYYU�`c`G�o��}LL�X��/��i�� ("��/cb�R����Vc1�<	�8a_��`�J���\�*���2-�+Lq� 伸�)�������hg ��C#���õ������7顧�#��DEE�C���VA?R�����m-�V1�nQ�z;`�L<�6������c�O0����$�]| ��T{�!݄MX�]=�^Bo�Ql~�u��;��dC���[�eX�{=�t�+r.�O�iO�@p��r�߰�%��sZ�����G��*/_w���}T���yŜ�2�Zn�����%��v���� Z~C^�ذ����EEZ��T�g�*��"�d�eC>�cw�*�L2�jO/�X�Z�V�UOǱn	���\�j����22���۳�Q�S�������8��-mm�����y-{׭z���� �-���d��c0�v׮}�k�T�)�X��1ؓ��ڣC��%d��lr��~�E�ԑ�&&I��/��9aƏ}���rpp�	SA����{�n�|h���$#=���ͷ�y�W�<xWd�� ��[���}��"�G�A�=��䵛.��L~��U���D�eFE�ǅr32�L`
c��WUI/.,Ȣ�o!�S�&��M���>�EA
�(էCX��A?�K��y�*�N?�֪+��b�����b�޸,��E�8^��o��Ȉ% ҇��s�!�
O��%��|���pQ���+cA�n1�49�R��硚?0��>���G���[Ž�r 5����3%-m|�|��Lk�a�CP���sd��0 9�M��)L1�����j�:�&�[ȶp���n�#.\���àʾ_θi,�BG"�^]�&����'(�@�8���%�e���H$��5�N�K=6f�S�M�2ޗ�Lغ �]p��N�G)���1�#��@�V�S==�nn+��8O�-v�zi��OU�Q<�[;69�8�8tC[;�r���)�y+a���zҗ��� %��<�}hi�RT|��	��!�"-}��_�&���}[t;'(8Ӳ�6�mf�VC��͛[�k2�fFׯ�O�rꆆq�y�!�V�%����,է����. ?�����K�sr���x�K���&�>���?ӈ�óS��h��	5��^����#R�B����{�j����=�4��$�������T;�ߺ=�	�|���'C��/��UTt�rs�glb���E��l���[�m�>���sbi�ug�,��2B14�p���xg6r�~[D	�T$4�"�U���G[�vTCb2�)2Ը��;O�4~����˾���?3�5뉯oG[[B1�K���m7������i*O76<����[�:/�t�O���/����G� �������"�8�HZ�2�%d��NsT�A�������� �Ї�3��\�դW�Ɂ/�ၐݍ�=� ��7��T�sɾ/�f�$<�
�`I��m-,,
@���������Gn��2jKR�Xn�y����7G��������%�߼�ˍ�Eo�m	�y��*�\,M!����\3�P3����t�����#�n�����m�)Jö��� 0223�EP�j��������/GJ��ѩ#�����#Q'Es$y.�:p��@N ���Ɏ���W���r�h���K�I�EPo ����544$�FJ�#��o:?�0��BS��9�JI�>�ϯ��t�,��X�&y�ц�)�6~ۏkV>�,�*.cT��	�-f�	�QI;�������S��
.c��xkb0�cc@gddHG��ە��ɞ��.���ʦN٧��>������>�100���%��V��t��Gu�I�XO�ͥ3���r4�0� ���p�3#o��������˥��k��"s �����!�+w��rv.&''�`p��L�	���m�\�_�����N-8���7���#�QY�Ϣ�3Н���u�N*���)��>�V��/�X]Ɍ�7@O�U}�����s7>��]��kT�a�[k�����?��=t@��b�yN��K/��E�\|8N&߰�����WA�s�ʅS33�z��e��������\>�(�33wlm�/�|��<���g2a����b;2�-'�V<f��<��_�R/�lV)bf�2�/�F�9�=���@���-�-���X8���7��$�p�|��A'�>��T/�s��Rl�4�9����g���U��'��Z/���sny�rH�路5��_�da9���k^%d���28)|����U7^n}i���/b�r<��j��AmY �wxa��a�)��E@��+*���1(��Z_M��lY龜���ѱ��3Mh-��������Ѷ�����ܪ*�vS��}]�zi���Dū�=z�&�=��*?�����*C�z)��*(���

bdb
��y�V��l<�����Q"�U d$�&{4��Ӯ�1E��wll�s�A��M]]�_o��t��lH9�Nw��k�kl�"���)�?|��ۿ�ee������o��iu���7l�v���d{k�2��_������ ���1?-3S	dU۵k�ȵN՚���^JJ�m�C{�Wf�R___�������i�9eאp
*?�|��͙�M�Az���xD���9�=r�̜��r)�}��k�{ȋ�� 7�݂��22��c}����5��!�3�6S�q����;wwP�W�<z�Ƙ�0H��O�H9�H�� ��R�-S\�U����ܦi8��A�~M�����l��h=�ѷ�%3.##�a8\�bq�c����oh�֌�r@P���+�qL����lĔ2{�#�W屪�Lݨ ����KnMJN�=,����eaq�\:G�zK�h�D%�]տ��<��V+����ϣ����j��X��o�@0���uk뜜������~��G�C0$=V������m:.yй��f������մp>oJ�)���27�?�w0Zt��"�eok�w�a͇�t��ɴu���ԛ[��]�)��n/�Q���"��X�\i�[��S!]��`v�n�(l~�HT|��u�I�K�f���s �,k��[�LU$�{�1�S�����J�H[���yj�UI��1�:Ձfj�[�E��ښ�6d�쫘�R=~���Y�NK�2r�Q�}�^�����Q�\��������z�o�Ń7��R22�V.WNg*��RE�`��l��=4���!�������+3�m�f"�m}� �W�#2��YYyS䩩��#B�[V�j�Z��u�ж#�B���CY��M�ϭ�rC�f�C��X���o ���_�{��n0����RN�xS�蹾�*�Bv�����8=��ud/5ӊ�;+"�o^@�l��szʤ�2.=�x*
c�w��a��;M/n�w�"��6������2�����$D���NEp��鱵�\�lm#�p�LvDS!Ō0pbx4%�����9�ct��L;t��5Pj����xT�:t�1�㏯ۍ�[+*$�DD�	xᆲ�O��@ H�ů6�ihjbєBUU�z������t�2�ʙ���'�5s&&���Z�)�,!qs�ȟA{m���8J`��.O�!����������7[���bd嶹إ�F/&*���BlK�ugJiߔYҋ�_��R��i�����A^���F�7�egV[���@ݥ��E�����Zfnn�uX����|kfR�p����c�����)ȫu�z�2��k���c�����N�����׃8���f���:z�^�|�Ҹi�������lK���p~q�9�ܸ/�q��
 ��Ue��w!_V���(������-�q=R{������RT˥���@��[er�b�ov_SR���V��8ͪ��\N��4)8��h
X��{0(@;B��ʝ&ú�������8��QQ��E6�*㬋���9*���S���� ����:��@޹��ϫd������01-MAf���8��;��KF^? ����>A��
˧9��{�<�s�淕m�HOoS�K�M����PF���?������rR�"�]=ř��T��W�o�h��"Vb��	�u�Ā��KF[[�����@�?�LU��oM3��F������x��S/k}[���~ ���<�`g��{�p�r鋥����N04Ȱ���6��k�p��҃a �;�Ǯ^v���ÅK��_g]�c�p���m|\�eLf��$�>I�B�R3�&^r���3u���H�B����8PZ��-��d��¿^o��R��tLM2���$�������aom}�Ǽ4oMOP�A��s30�0|�M��ltĻѱa�S�v�$R?2���ܻu:��ނ=CO%/�Ï��x������(�E*×��j���9QQS��GB�&{�3���@�ݼv͟���x+���^C����*4�<�:�\��zV@@�ҥd��=E�ҖٚAl�}��Ǘ!����&�6������)5��D��z�Ԧ�� �z�2W�.&���#,Z�x5������i�X�+�齖�����nnn���Ծ��Y�>@��ȝȯ�=XXXX����\�����(����qm�\SK뇨}H�{�nFF�v0��3��d8�i�?�e~�|����)��#���s�L�<����SR�������P;y��W�G�I�s>��	�me������T_yG{{"��;{�/nȇ��m�cDbmX��;�4�_	��+�/ ,��*#5>���b�Q�ƚ�dK�7��3���"+��ׯ����l�u�x�G<n	�^��c� !!�Aj%���#_�G��B�R�{��bsTA��ȪG�G��2�^hW���X��bp�fP�4�����O��w���\�D��ٳgL,�����ee)K8M��̼>p��m�yA'����!��R_.
߮aVO��s����:��|��X�N��䛫Q-5���ʥ�{���5�g�7�;�<ڋ�r!�?�<�3�&i�V��侗��C����bm-�t��#�W${��b��=�-`����h� ��w�C�Wn�R�QSN�8�����;��k�����:9�\�p	ԥC������Z����ZWu���+2S��Ԕ��ʀ?B� ���ο��1j��&���_V-3�4��}դ\Ģ@��"��q��6Tn��V= mXX���Ǩ��v���'��K�]Q�{��=�4�7���za�ً��������i2��d$$0҅$p�1$Z�"������]`Ё��I�< [��2ɻ���.�f�� 퇼�1> �.��ˋ�!±�5�5���^t��4?ww���P��p��߮��Y*�˒r{�gϞ�Xڈ�����KG<��lAӥ�B��x�GYGX^C��������N]��m8�cp�)�/*Ϯz ��{ [�>��--�T0�h��B�e�}��c���z��������h�)��4UT��,.^�I�����D!Eb��ʅRՏ`���Ĺ��:�b�\D��Z���d�~*?����,�v�߸d�~4��; �w�rt�)�������ݏ.��N8�Ѓ#�}p�j>~��{�-sW�����e�ݙ}�ȹ�>`���2���?T ��e=�hC�M��x�߾FY�\P������S�u�mq� @ �ؖ(��%8��?X�L���7��6��QkCX�\b�����)�sc>{hi)����Q�1,�y��]����\ۜ�ν�G��gb�ē[�Hŧ��/^�����&mȇH��Y@~r�;I������<�aa��#�x����9�8r.,5���d\��߻9vC��M�����=�1cff�d��^P�N~|�.���󂢢1�*\I)�L{��q�-Pn� �x���&�Eu��GI[����.�������G���T �W/_�c���.i gb`���cv����>:y�F�k�H!��{=Us�%���!=޵��
��o��~�1SNC�O �ssSS3d��/~�O��R�O͌6Eﾺ��vU������# �h���|��ojkG �7��[�����L�yI5:����9��`�j����\YZ�J{DU2@���Ƃ��7Z�?��!�zA�_�6�an������A.,ĪWU��4�^7mS���ϨJ��*Z��_ͱ� �j_�S����
��z�������?��;����P��E�a�$��2ʎ̌"	�D��̆����=��(YeG!+��9z����������s^������I�5�5x��5����r��[!s�冁>�V�63Q2��|�Yr4��^^�GM���	��Φ��z����sr�J/����pC6�W��5�Ё���MM� o�+.>u���e��y��wX����]9V|R=� <����g�� �!w����g` o��刐B��w]!uk�jp��oZ[����43t>���s|�=	l
ѓX�����:Y�w`n	8� P���YO21��NMJJ�y#������m`?�		զ��L�+Z߃�s��?�|ś+��`=�
�GW�&։��dGGG���������
@����=����[{��p���!�?� ���n���g/)�v��x3�`c3�$��]���t�>�q�<�450��!�т��1��v/!B����Y��,�;�69�.�%0��6XՌ������w���%&~`��A���`�>Ì2�7�Տ�s���/?���
N^�0��!}3��hY�=�W7�(��Dc���!}�il���mJv_u�pO�6޼2Gr���Ó5,m�saJ_��v���ã����}o	nߊ:�9�����V�.�籩n�c��9V�Vg2KW�i��g���!�!;���sp�9�a%�a
�92��HH�d���8G���`}��J>ǭeC�棭��Y&��i	k�vnIK@?�?�:�{��<31��?�ON>	J�E(��:�/�dZFo�\@@@ҋ���=��*f��g�o�;��9�U��/�Bp�N̩ʪ�/tI&��j(;����{�=�D�<x��ojz���K�� #�h-[l����n0S�I����l�FF�-��\<<��TG�[�t]�_�+���P��˷03���Vn*#�@�H5B�3D����9gl�!�xw�FbB�'�A�y����Jf��Q��#��~���榩�Q�@�.Us��f�_��%C�ˈ�@����w���'l��/����{t����tr^޼{�z��Ğ-g���[BAAA尣$k�d[�n6��...~)}5��)�ޝjb��p�;�c���A��@�iI5�Z���󃝷p>3�A%h|�F[2
�p#-���d�m�{�7� �e)]�iN�ݩ�N�۱���h�#G��^a��j�|1'''Y�o�v��>�V��?2<,Cz�����	b$]��E��-�$��-x��	|���M{�"z~~~��?�����[!����8JJʆ��1]X�e-y�{^~�޷�9����W1Y>�>�"�N��na�/�S4`�۠Z�nŌ�����H��׷x
f�����^��=��ۜ5�ޣq����]N�QQʉw�~gY=hη�����OCb=�A��OxNqF�v!w������+���׫O@���ѩg��'T����;���'l��">�������x���>��IX���C�.�Q�߀������)��.��y5�%����V�G3n)TEL߁P� �4�!;Lkm+/��V9���P��D�X�;#R^�]��.����ݽK����r2ekooL_�AM���p���SQY4%([\��Cz������I�JGʣ?�;���C�zܾe6ٯ./$k�l:LC��8]��n``��p�6b<予��M���߯�
�������������U=4=\�4�7l��i�����M����$����RtX�[��3a�f�/��IH?�T��X�ܹ���L��ED���L�o����*�3^<gh}�|�Ζ�Q�����0wt<!���0���Y,.A
���:9��^�%ъ-��Ba�W)սoWx���N��e�����mKe�6�"5 �A~��`�>J�����fiZ<jĳo�[��D�{���b?B�d��[�P 8�}�yS1�qHE�Ň���.ΎƠ���w
��l8���.@�t�Ê{@f�Q���M �NXw&�=BB~H�n��L��.�<�(Y��}]���������#����B5��x`ÂC]�,���"��5���X�.�o�?��Z�����N����,Y�| ����ҿ�c­�x{�hu8�F������qZJ��ݱW>F<H�j��G�7��������r0������L�b,���)ȡp��=��Uzª�2���Yľv`���t y��=�fE��ˢd�$ֹ�NX7$oڝi}��Ǝ�#2���$0���T���U��ؾ���˗S�����B�U�M��纼�V � Z���b=��t࿷��~�#��OR6��pSme��/�o6y�2ị����.MWW��r�UǶpn����e�UÎ���|�gk��ᱷ�^6^K��3��z�=�<�U����nM��������$ ;��%�"��3��zo� [��Ħ���o�t45[���k�Ӫ��?ZU�٩op��)x�\G�U�xE_�k���P���|��L�g���E��
`�[�h*!�֫�o�!~��ٯG�僝�A�uÜ�_�6����H��/rG6k"�2�a���`�xh�@�i"'/�ִn�����.���V�s�q$h������.���Ox��E<� J�zY�ʂ8�Ո�T)k|	����JQa�[�z�)����I�[K���H���0�!����,�I�b��\Q� ���Mmmȍ&��7��X�cu�6�[#��b��x���G%�>��h[��^�S�7��������glVg�.�3� a��]A=���0�� 1�{�r��#opn�ime.5>��	�� �z�R~�EB�HJjƱ�K���s��"9H����#ddd(��}����_�§�&��>�a�6�0��ɡ�@����g��^cq�ca��r^��M��I���S��k�\Z���䳟��g�����J����p�{m��:+�#�uc-]�*�O>~�uy�&ș�m�vپz���������~G�Hp�l��j7����cGVg����K6}a�/�3�:��CN|�$�K%zs�;�����L���)�^�;~�DB{ayy9���Q���*^�'�Z�w���oV\�&FG��4]`�LZR4�󂌳�U�V� �����������W��ƖPʗ`ϙCC��?>����{��AU�{k%g���F�9[WgL/B>ѽP͘�G>�v��]��aK��%)i��742:����}��lN�jwJ�B3e���G6 +�KBezΦ�{bQG���!u3[�ق'XM{�$����y�-�-�b.���[;4�0�m;��6H����D�6��kr�dׄ�0<�%Vr�]�Ε^1�(GH��J�w�N����\�Oc�l���N��g`x29������O�ioOTt��o�`W[6w���k���V���43|�mN֘�X[)�SO$h~���e�{�''V�J�I2�겉�Y 
ѠFk�F�1*g��������i]������TA��ec�{��Ivo��L�������,��S�^�����%�ZAX��Azǫ�dw����ɾ�d���6�^��r�=��KB�KL����\/&s����O�1��K����&JcEɒ��c�)�u�$���P	 ����ggg,X�?��k�om���TX@��U�S"��#a�yG�=w�\��hĵ�+^����cY��2ywDy��r�K���Ah��ԩ��)))��
/e�{�Bb���XG���2<Wr��'9�pŘs��
ulO��0�4�<��ٺ��ƴ�n������x��${�gY�+��J�l%��6/�U��ʤݿo3���I���صe��+�l�V�����e�&'��5���Y����Z@�C}޹�O�F������锐��7v�t1Up5��٩g;1�@�����(ڽ� �6�̰�(5���p�$
l~	���>����Gh�_(����߷/��{�$(ꐓ[S�|�r�~�2.�x��"�~�|Zuu�|%[���ڤ�jV|�G�>��������'�k����*ǐ4���^�&���qcgg�h��ť%�e�0�X�'��FG����	�c���-6��_k$�߇�~vzr��K���HA���d�Ƒۃʯ_u���N�|"�9i7_��Sorsz9!yO6k����sj��@�.�9%�GL��.;X��s��N"�&�|�#��ɅO^�~U�#�qAXAquFu��_'=k�~�����;�^��:	�,�u���v�#��t�nz��K?s�t�}��sV��h_����em��扠���ϗ�~+Ks�)*���!�^BC�n+��Aߴ�:�n�xqzuu������(��U}�1i �wI�1���A�C���z�,:r9]��Ҙ�l�6ΟP�Kx	���I�Fb��e&V�'��2��<�L�؜��ҕ�0teQ�+}�F�RY�iHJ�k,�[RS�{��1�H[Z�Յ!�b%�+>�Q�����D7���b������������߿1*���nBF���8Q�x,�s"�.=zܒ|��޸�������f|�$p>QQQ���8�$�z�"<j�ؑ�J�]H������ds��"!5&��|�q>e�%�R��ߛbWG6e��T;B�����
����Jf^��f�(Ő��Ӿ/�P����^��|�����f�Cf�o������eH'�*΅��k���x�?Yp�8��o�zVƝ�5�٢�>��S�������#9�x-�_H\�����m�ݟ?����;_�;�Y׵9X� ����¶k/��0 u���z[s���9�8|�؋�a���E-'g��E�5'�2!�h�(�?⿇�X
�IN�T�D�}���4{s�z|���qFB�	��p������G�&�z,��_�nJ�г�5���\YI���_w�}l��\β�����UD+�ɬ!�lL9_s�89ٜ���d�o^��Y�FX�g<r:c���=� F/놱&�Artn�sŋt�z�%KX���UިX$�E�.����Ob����/q Ru��%�:.�q�t��!���	�I::j��k_s?��=w}s��N������k�+Yf������fzu��m0W>�k1n}u�!��woy3�L%����Q	�椥C�׏A&,]L�������L�=��T�u���Ȧ��[ޙc�8����j��ſ�����2�Kޘ����p`��A��߶��a��}SC�i� �N���9��c?�.�<|H�S�n���CQ����^���v�;a��1� �ef&j[X�<s,���,���~jk��T��&Sys���I���|���)�y���G:��~nś��)���f��߿�@��G�7�|��(�Zx,��8'L�Vq�קUn^�����<�E"�MCD���Ov�9�=�Ì>�^V��_Ǳ2�9@��������]U,��2<��k5�32*��ux�
7E�RR�nnn�(<b^��E��m#���L|�� ���ְd�Ùi��f�ϟ��U{~�a�5��%�TwpR{N��Z��������!�d�9�u����_l*S����Δ3���%M+!!�,8b(a=�P��(EƜ���r�k�:�ҡ���KW��C6��{}����<;����9�t*K�<��>, �<��7��j`�B�`fȾ�������kM�ݝ�����LCC��t[���u�e��ȸ]h@��2J�
r�'iK��!�P���T��c��RA+�bW�p�op��ln��X/I�SG�����sbC������}���C��ȅ\x�¢�ۨN����W���-?��'�s
x����,��3��ɟI�����7�ە�o��oÊO��;	�:Y:�ts�j6 ��M�Fiz���9s��ǝ^�Ȝ���=���!��.?ʃ�	��ŵ�4nu�~��M2|�䯵��T�`W�Gw��im__��1�$��Wk���;��l�33�Ή�L~~����C!٭7I�&�k����b��q�~˿F�3��v- ��E{*�+K��;<}0q/�(	���;�4v�;�/�S��Z�7'�ixHA��_���������Ѡ��� ���͍�\����es��F�gߡlX��(�P_��k7�4�ⶳ;����Sr�Z���T����V1��뫴Rk��A|�ccR���/��F(++?����),_�@c��q���V4���n{�׳���'�}���f:i��c���4V��[��tȾI�H	�'n��-����H`F����O��geMj�T���{����y�GL�À�ƞN�[����b�@��٘	w6'R鳘֞J���	dd����egff .ٓ'<�
Ѯ�RѢ��
�b�Y�v,7��w�n$�.�a r����Ԗ�b������~O�>u���
�f��h�)�2�]_�qT�Yh�D�t67;���K�v�U�^}���d�W �;2�;�V]>k��4*ֳ伋0�·�+�E�$�������6;m�B��s����������U�;�ɫ��o����PEY��UW�[!�=7�|�d1���糁�a]m�G�ȥ���-���lX'�a�z���lRY��N���"�8~���tc����	��ɘ?�Gl͎R.���q9 ((�"���{�_!�=�ZGn�x�v���Revf�2ʦ�(Y�599���U;\�ϧ�_����)�Q`��$[� �@�vb��C۳OӼt��u�<�q+��:�R��qi��˽Rg6�t��s��*cx?]�E��y=�e�ȸK�v�
�(\�mxc����?o0���_���\�.,Řg����M���������TὮ{xxL.�f�)�^��v��}z������ 1ba�r�6=�{ϓ�9'�~j�_ȿ�%�����z��ݡ�1��}���<����`��!���>���ec{���0�l-mA��n�=SFr�9b+G �j� ���a��%�>o8d�h;�u&|x��eMĉ���Xamd������u���L^s+�x �d�o^�b�i�q%��O�%3���H�>&���J1j��,�gR^��ۀ9oQ�������́�Ͼ�]�v:e��h���TT�ͦd�<�ǚ����*�Νkx�+ 0[ ��Qnd�gzr_�&�'|\;~�^�e���ɺ�S��#֦�k�U���<�򓼜���yx��؇��I��R�J��z�1��!P*�;1���Ǐ�p�(ö,�'!^166����]o��F��o�w�T���MV�,��n��d�L����(/�r�벫2������j���]fɢ���BҖŁ��_�G[Ӊ�g��UV�݉�Y����bQ=;?T��X��^p�D$x��6�X�sK����y7���!r\s�I��22,�Y8�;�U�����ɚ�L�5/v!2猇����t�]5���}}u��T����)���r���}٢9ˤ�o=�rʅ�N��9�?Q���J6w��\�=4k�sJ9B��̋g�Cm<�M��Y��s��A��Q�޶*�E�@{^�^���?z@�E�3�;�lg�j����
wH�	곩�#|G���оwρ���ⶭ��y���#��Dl4�J�Bt��.�>Y�1�Q@;��Ȯ:���!@�}}Ey}�2
�ǅ���$X��i�9JBn���g|��!����>sN��ke�y+�.97W�x�_��q������R��u��eA6�Kk�Z$ӿ��f�+�o�iP����7z�)����J��s�Rb}|4�VN޽���|�X��S�4J���]�0�X�J6���K'�c�%m7��Cp{���!�a㱯Y�7R���
���Q�
v󿿃g���Up�z-�m��ǰ�.r���DG��?BC�X]S�1t�vNN䝪���B�1�_7���b�L�n|����[ 4�[M5� �3Ҭ��"\���e��֝���0Z�{�xW�^���	�ί�m����d:�\@	�(���/W���dҸg�}� ����h��Ï	�***B0�n�:kW����a/�f� ���(�v��fV�9'<^0��S�y%�a���e;�q�>g��ӽ*�@U���*�}�)>�^�$1'C���v����|R'�E��_l�t���HOO9F���u4^��ӌ>C�=X����1�`��t�y���;;� ��Ա����Y��}�Q4� ��R�]���A�p�X!�hĪ����n���$k������.��/\�RC>���)�L}t|<���濮0��I�)��0������U��O����i&��f+z���eO���Vd1�i-lI�NTI�7���P\,	�/CR{INN�7?����Al���3�N�� �R>jۖ�pf}�-�������U͝SAZ�K�ri'���tT������J�Ml�#c�=A�u��t���s���,���,��
���s�����k銹�	BS
�jM���(��і�yNXM2.���o٦����O>�{�/��UFگ��1�:�����x?oi�pt���K�6/gBn��Fk�<&pK� �F0�yp�	�����<<e�YV��J@FH?��le��K&%E�����ɿ�� r�]C��|H|z�,Dy���`����r~���M��ɗ�(V�L���	�k�+�Ʊ�&�Nɚ�`�=��22����;<s;�h��lj�/_�D!�{����"$�cT�ǡ��>��'�{z��1���X�z�>��9{��L�V语`:�YƲ#�l�B{67`m�����~��q�t}��;E�{�|�兩�Ǔe dkA��),T��q��Q,٦u�l�w��P!$Y���M�S��K	pc����D�!�l��To�%�C}�
��w�ܲ�Y����K���R�ɋԽ7�vn̪�ؐ�Ǎ掻_�$�]ifAO�!���@��o� �Ìt$VV1�W9��4�m||<擖i�3�CY���=��.�Q�N�`����������u��ѣ��e+��dee1�%o����\�(B�Le$ ����nAӌ�)I��wpE�������2Ӻ0��Q�ds��3=�p�4[ces�i&9��Z��T����7l$��@��zgtb"����P��d�0>���Ϯq���eE3I�!�V
ԙ5�N�>���� ���	��L���g�������c�ӳ�9��ܩ��_��d���|h�[dp$���d��(cə���l�v�켿��^�<���cfz��V�L?�(�ja3M3��A���W`��B@�;��|d��>/@=�r��Xt��j(���6���+e�ِ�l�����������X��z~����z�5H#$�5���V��2�s��N��)��2U���/Vm[>	�H�+m,�w	�\��u��i������Ӯ]����� �:[%���ɻ-��J�E�c��  �3��q���h%4��Z�BfwF����`���jF�/��h)�4o�+/+�)r�����ɩ
0 ��,���]� ������J�ׯ:���!FÚ��;��޽;|-W�]I�_mm5��y^�KH��n�0�.���
h�<1>9�c�!Fl@UCC������1��������[a@\���5�b׎)͟w��dp��/ ��H�{!Ι^�� g�za���[�H��	��@�>|��)  �����!��?�:�G�+e�S`=\��*��oG_�������q�<�eH����W�Q��Ҁ�������@_^�-����Hm�e�#�8?F���:|43fn������:t����7>z�Z0�h�g�C����*ze>{�}�kq~��=�:;A���8�4vv259���d�p��c���*v��6,qR��s��Y�2�����xK�}ȋ�X{4���T�IU�u��V�- ��H�<ۃ�&W���//�N�ܺuK@\��×�*��؁M�����]���d ��0M�7W�u�D��6>��84�6k��`�ê������/������%g&Mh&��Ο�i�>A=�۩��mll 9DbYܿ7�w�p>�(��
~	�_�ƋS|3��M���KJJ֞����U��5���d�Gx������b�kf���������� �N�J���y�a�J�z���.�R������o�
9Q�R�N�ji��T,�L�5��������4k��"4v���RѤ�ё,@�Gs\�0^��9�`���1���3/:��lۛ ���o�]S�x�I��1ͤ���F��%Y�LP�O"c�y���'�4�����_����hu�ن�UTD�K]�=�?u9��9#�n������������S�Q ��9�,� �@�HK�En7i����z��P��F��_��^���x���ܙ3�i<�W�u�[6����6{�亗q���o� ,�Sz������T�6l�]H�n�S]	}�0I�T��w\ٗ+��:}f�Pe���鈺��<ɱ� IH�ɵᖦ�LJ�qP'2�6�TϮ�8�*꼪�]����X�:n��y�?��vcu},� !c1/��P�o�I%�e�����]57��R1|_1�&�!�q�K����s�X�D�-D94:|�X;���Ӗ���@NR�*hA�����V����˗5�X<鱟� �
�w�n��'0(ӓ���%<��jQ|����T,��L��:�֓�6���f���4,�����g]5�q��x~��e���f:��p��^��y�.�*-
;�Htǈz�N DvD%)����bX������,������-W�^�ttX��RVVF�M��%kܬ�X�%�ù�d�z�+�b����ъ=d ���%�b��@-��_PX�۴D��Ĥ�Y_>�Pcω7���U�K%����o߶\����M��:ye������vN�<� ��}4Rg�N�	ؚQ���C^�
T߇����ﾻ�M#��F���ۋ������Q6�+Eo]�eƌ�YC�U+����ommEB^�G�<�Ǉ�Tp{Vyy9����b��K�*[u&��aܛ�K��?��+��8A���E��'&�a�#l��j@W�	�����3�`�����:ŮN�`2�p�Y����4�tw�X�gi)W��=�aո�v�sn��sY!��_u�1HZ?�"�o��N]]]ķ��k&�L�B111566���@�m��eW�vf��������Vx�ˎ[�\�޾Դ�*�ܗ',S)����D�v;�xZMG5�d�BAn�[��_�+�DMu�`OC��2Ey��&q�J��!�S��d�J�^$}��&��Mڍ��d��|�4}ܷ�B!�o�U|���1�z�w����wZ����:4(ص���/^�jki2;Ғ�_'��R��KH�)�DM���\e�P�4S��t_��$eL	�l��bH��6���-�����MW�#��t�3��8��Z[���0�;i���b`�,c��u(���)+��Բ�h�"%\���7�]�1}^x�<Rg��I\���5OG`T��5��4jv@K�9�A3�OO%�>W��ف��iI5�*p"��'�2&��-q3�������?i�X������#35�L���T�셠� 6�'`�7�%���F�b�4���sqz:�sfL|Ȭl�E'R�K?Q�tI�ӗY��;߳�Y�к�%��U�Q�A�\���v�jbbb�V �Jn�Px�拧5��m��?�&R��x���]�ǜ���È���ӻ�AG��5��k�"v��*�Y=<��e��0&�"�����s�w6�}PWA�v���ںg�5�_3U+� ���E�ˆY7~��@t�z>��~"��
�R|� *fʶhs���	����P���l��5��ߠ0�=���N��ۍWg�Up��7	��=K�<�es�G�uY;���{z�nhbӯ�:|��duuu�~�.9�
;��|yĉ��x`�L �FFF��I+x����V~k>x^��9.Mܜ��6js�˗�H1�[BU���N��c�R�R��+r������o|���.�K:��v��*NP>�`�d��=��e�'|?+XV/���)**�hS6�"��199��F�D��]��=q��N4?С�H�ޑ��4�7���##�\�o;D� �:pVP��˗���`<���}�@�$4��k����+�m����WݘV']o|R��� +��Vf_�Cɧ��ǥuo�Pc�%��!�`�M`iRNT�R5vZ�Yƞk󵪞��A8l�r�s ��FߴW�����Bޯ�@_�ћ#�h��#�7D�IA�cL<��9o��JP!�%����WZ��L�m���`���_�8�Nd;������l���9��"֓���P!��#����n��*`��l$�Q��_�ie�3D���[�(��"��R�fa��%�s��JL����_�de	 �7 �9����8�x������	o1���ǣ�P.����(��e��7��<��Mc�
}�C��N��H��Kq��6>��^C���< F���%}�%����=�N�t3�V"����?��v�cUEfyڗ�ճE�HR�M?����޽{�L��ƈ��d�ƺa����2�x���U�]��<����0��K�osh�V&���K:�\L���5?y�2Q<�w�[Z��%i)�%���/|�"6�����ox�KXw�r!O���A	����ۨ��<q�	�Y�ѭޜ�N��s��	K)!�]�.:����9xU��;|��7Y�vӬiȈ|���I��E�G@�H�B����# oL6�đ#��`SLgS<�E�A��45��Hn��wm{'i2���J��`���=u�
#��☸8�����$3,t�����/�]�I'{oQW������cŐ�C$!�@�W��� �*�+t���dl�q�X!䑑:i(�)L�x,�$68y�`��N�<>���1�l��X]x���ĆG��\)�Jq�l@6j@�_�QQ& ��ȥ�/@r�`�1��q�?�֍�� pei�fue)0["G	���k6���[�0l�f��Kr��}Y�.\v��v���{ �B��r%�����El���i���~,tP�8��W�\`H9�_c�
"r�=<
1��_6�|�r1��@p #ؓ�	�pT�~	0ߨ�-bnQPW�c�sil�8�)6��+�ڿ��p�M1�6/�5N�M-8h�"�����DX�)En�CFpN���î�b��;����5�4<B=�/�lb��;zs��8k;�sA�--�����рe��zy�9�TW��X���à��w�	�DC�M�3m��p��	��8t�^#�S��L�� ��b�R�v�yk����|��C����rB��6&�1�Ro�2BU��]q3�v�
�W���(���m//.�e�L�'�0Gd���?a[��C�DϿHIdaG)��`��<x'7}�*Oя'6,��L1�mJW��)41��^B6Û�_K<�ħ��r�
��%�74��<u���ɲW~�G��� ���
����d�o�y��N� ��x�d�I��$�D�m3
ƞ�x��XI6)��cW����6s��`��v�9[��S�Υ�F1x+�� t���Ŧ���qt'05*&777��]A-ň� ?>���F>���P!�D�ut꽨��d�$��в���7�زI����6Ƹdx�����1*T����q�t^]�g�QRT������������k��4v�N[B�1��܁��=#'Ji�S��Z�����7a�	�{y�}�/~a���`v��UMT1��>"@O�Uv�M��3���ʘ�d`U�� ^1������]���<�2͠���Lc��:��G�&eg���;�f.[���-��ê�>����}% 	�-�
��9^�3jFlc��P�DD�8r�Q�aU��m���R�����wH[C�z^�����{`�m�ݢ婺,��?�&�ؕ�J��Ρ��=ֵ_|]�Y�'R=��:�F��:q�,�D��`�M5�Cu��eN��[b�X�n#�W��{z��~[�/A�7'��c���*ߛ�����Ӊ��[�Ꚛ���n?X<�FĶ�G�^`{�8?!aay��B�t2GͶN��fMudg��؃Jԣ �/�'y�]u���K��L f�����2*�|�>U��C��Zhb�v�4Ϻs�Z߫���Fvr>��?�r�@*������D�������|����s�!��\ >ĥo+�Y��X ���4`|D�#K���r��[��)��#�|xiݵo;0}x����E�*E�Q��[N�_>����&kX��,[�ͣ�����O��;+�b�ص.�"e���&�����%H���F؅
���A^�o����sL�E�ޕ��ʳ�������r/���r��_�3:�8]46f�3�5�7F(3E^�"��c������cm	*D���*��e~z!z�����, V!�&.���w�b��N�(�zh�km�8�ǫ zv@���
�w�w�Xێ� _�C}Ұ>��>>be����;�-�"޵"#�'9��(�����\��LX �'\�)����o�EK��@ ��b��s�(�#�(R�?x�7ik�9����>��CI�q��YI�����Eٔ0����Q�T�|��H�`��V |���U&��hh�`Z�!ݪ�:p�	�oT�����58_$�6�6%W6����{�k�_lT�зb0��_��+"	�:v��� ��:c1=X����l߲M��;Ը������������  ��q<hr��/�W�:և��o��x��<���2���4oU���t�Y>��)�ڠow�9u��9}�`��nXUc��IMScOO�(!�4uL�x%/��t3�L�%��	2Q�O[!K�?q�L���ZPm�hieeeT�LLL�������4f�
	aDrlw73~҆w����$�y �>�1�6X}}up���f�<�h}t�N@��$�r%n��.�c�P<y4*��2�b��J��t�pD��y.��b ڮԛ@�C�ǆ���SZ��M�#��⣸�#�\Y�M�  jW"�ş�~���Ëy���5ӈ^Y�ĉ0��Y;?F��>buU��vr�����1
f_rdս��b �A��%%%�w��[~kr2�KY*n����~���AT���!�j��V�.9�7?�g�.��&m��Hǥ���B���5j���(��9�	�?��t�)�0b��+��6�I�r�"�2����-�; >���<5jI��$�(�S�V,P ��I����Ε���]�ג�I����Q�!z������`q����R$�A����{���B����Í<O�d�mmm��fre�K���\�#�R�q� �����k��*#o__y������\���Ύ�u�����c蝘��O�G�|분��];w�{���[\vށ�v�o��]��%�����4��0�|s'�=��?�pǼ��Ai�W!<�=��=4'j�.����61��d��������O+��o����Ka	�t�
��v���b<�ũv�H��k�%�Ԏ��^8���"�:�̈́SX3���MQ����D7��l'�<u�Z���Y	� ۡC�$��X���t���@h%%%�&j��s�إ���m�����.�\$�wqǾ�g�&�2H��p��(i�-1��mf�<I��{�1�>w�c)���ҵ������ny��|7[�z����9֯U�*�f�S�7n���q>ybC <�ã|���V�T�K�X�k��ȣ�w�q���=�o���ܟ$�'s��9{�\[�A� ���Wv�z�N���b�¼zO�K&��n"A�L��w�|��7)�m�44��J;g�Q�=j.AA�Cr>�V!�u���Q	�(��N����v���<��6o^?'oٖ}���@S��	��K�Q�)Y\t���Q��3���eH�<�E���'G�z-!�m��ޖ5mJq�v�L�9;�ggg��&8\Y]mQ�M��j�(��,c.��R`;���`�-�D����֋���񥩩st;a�V�]�D�����*]�"����љ�G�cS�K3�Z����AZ���7o��47�`�ܾ�d>��g�����l,�۱c�߾}ke ���}��C0��O+���$�B���%���.6'�k�*�59=�ei�4��S{��T��DJ2��<;��f[k�8J��X����M�]^2��(��[id;��l8A��QUUe���A4���y�<axWFHO��P���
�5��I9lz�
�ѣհ�7�E�S����|]�s�Ǐ�A��\�8e��O݆�7 ���!j���'���i�뽤�ZV۱cG+�[�^�X���161Q>��l}��]d΄�99��6~��3[�n��@r������Ƞ۲if81vĹt)FAAa��e-yJ�	���o����8��Gj����Mu� 'R¦�ALb���k�s�<>����d�	�
�ٖ�Nvv5Oϒ�X)��ʄ!>���cF�V�;--J��,.^28{Ue%��g!��"�L'�x
^��l�XY���F.ƚ(X�KFz�����~����W���}}}�/��	��yt䈞|�&�S;4m>��;�_̟�]!�����{s�۱����\�b�+�$ua<MY&5��\7 �66�{��;����-�W� ��}yk���Q�3,��ʨ���P$�9�j/�a3�S�:���Ѱ1�K F:�_Co�;�$����ϭ�xyj��}��T�j�� <<�<�Q���A�m{�H�|��ٳ�׿��-\S�`7aUEO/Һ`�(��U�b���� �M�����s�����=cqP����͛7cB0���)G����Q�#H?�nt���]�`؞@�-�=����U"�cE����qZ����k���q�ϔX{)++��G����ꏎ	
B0��_���:�������W��W~�����ã�$1H�2i��>!�����I<���6
i=Fv�U}z�n�v�~K��(᫥A��6�%��y`�M��l�J���ƺO���9���ʓ�iC���
�lA>��-���/vc��~Z����Gg��f�����VW���M�k��|����Hwq�����v����ߛ�@Cn�5"��	s.p~�D^�+���0�)Q�B"�����A�?� ̥���A7ְx�qig!�L ��ڗ		z��j�����6ň�G�F����KD�f��<���Zъ�X��'�f)�/y��b"�i%!�6g��"��3��Fo �T05}��@��
B�����Y��M�B�Xu�XX�$�a�6p�As]������G�c/]�7�̭$���K��8f�KW� (G̺�j�SK٦uX-�8ڦ'��?g�~�f���%�/�m�f��� P���U��C�g����?�VϢ��0�킧�_�^��|�g���.,,`nFtƝ�1bس"#1Jz[���] �7�����=/�[��Ԃ�p��6~��_Kb��+���rJ'��
������DNy�2��S0�Ϗr�:��]��!U�ܥ��������c_A7Gni�Ku���yA�5h�96B'Whllf��♿p���GˇP��A�W]�enZ��˿�f)���tJ4!��K�<GZ�˺�8�W�{_�iQ<}��m�#��\�з���~�q�^BX8�%1���us��3����X_̉�Vy�>��v�F:�E N��"�U0��tI�>���gG�R�⤵3�lC�>9)	�5\k?oG.��3wy�u9v�Xs������ȼ^?12�p��?��y98������߸����$����I��s����ꆆO!M\^�0M��'Μy�@�֪:���`�<���R�����,*o@�S*ZZa_�|I�Uh�!p��5<�c(�6�4O7(Ԃ�E����F��p�p��ni����w���q8}้��D��x�n݊E�����}x��1H�=Yc��D��W-� ���P*�s<�V�/�f{�W}mw�"@�7~�����۬��~w��h%�����]깂oR�m���3H�n�D�^�Q855�8�'K3���a���\�������!W�#%x���}x��f}���n���� �=�� ����Hs���`{S >���uJ����"DKy���	��k�x-g-{�c��)����-�Z�b�b��]���q[\�V�ܮ�n��B��D
"f��)@GB���t��f�]$��xg2h��Qϛ�>5�u[�K\>���e_�in\��եtA��7��0�|���)�qV!!���������U:h�8�� I�9������Ш�T�3OE�7m{.N�����o�d������g���u��h���H#���|�����x0�eV�H-�r���Ҟ�w�N��			m$��@����u"y:=<<鿥�k|{�A �[��f	׫�����X����=z}��9�K6��W�2S�q�.���4�<�`Q��Xtc�u�]�����pla�^�@Ɠ_��|}wgMy���p>#��}��׃��_KS���;���	+|B�6HX�L��ʮ�:٨��a��׷װ�Ѱ�^��܃������������C�����eG�������ѩ���ޥf� �m�)f\ �����&�Ϋ�y�(ʨ��\:x�.��	�{3�R7o���S=1���6S50�!:��>�h�gu᣿�W�r�?&x8���m ���o�|����+���
��~����b%�
� 9���䆿��o"!������Ν;SK+�oq1xC�q�G89����v���禳��[��y��}����������/^�@�?/+{�Hp>e�9gg��a=���:T���ޢ���m@����e֛������*�/Wu��:L�a-.��@� �U�6�gq��+bzm� ��膵n��	�0�C	~X��!� ��2�v�9T�L������ �9�kL�ϕG�
s��D_�!9��Eg돕5��4�M$��}����XI)�rW�3Ĥ�QY��Y5�&��΀E�tH���)�Ǥ~}qn"��� e�S.�X�����{�,�.��	���܎�n�^��H!�99���Ь�l��� ��oTc3$=�E�8�g��s��gJ�����rRPx��6\i2��Dl<��������F���~�>�˹�$�Y�b�<���D��#�%�f3ed�8>���dsf�R�zн�ebJO|������-���B����ݯP�Nt���	˜�o��	j$�",��d}y V]����Ӭ�(���GEM�J�dx�P�9Bh$B��$IH�M��T2���1��)ӷ��������>�s��Z׺���9�]oa0�����΃o޼µD	�Lۇ��؀��ud.�9��6q�Y�f���]r�"���Lj��]�.���ǀS��˃�!=+ˬ�"��W��VLq��6GGGC&�0�l��	o������H�Ͳ�6j7�iP�*0V�YV����	��}�e�f)K|�f?ծ�e�����j��M�����VVVx���DK����8�A"egM����B'���d[�9c��h���y��9�Z3j�PEL��,3��k�.�
̿(��n0Z�o�\�S�5�w�=)-4��&��o��_s�,����	��>n��)�C��yC���`�A�=���H8�Zz*TG0ƣ�M��< �Ͽطo37M�w�}r�_Kx��6'�Ǘ|}K	xG��VX��A��n4�vd��9]�m�U��r�:,��g�A1R#�̻�1� �i�)�#t�;ﲥK���,�3��ؽ ��bdKg8���R'��$K[�w��9
r�r���el+T^�F_I|�=x0� �+NK�sO�'A��O����@�ƿ���뉣9��p1�{�e�W{1I�O@�U�.�!߿O��?�o^���O�ff*Q 4]���{W��)`+��ݻ�����ծ�Qoe��_���20�tc�c��s3���C������	U#v�ͬ�<~ϩS���@ӨV BWSq��8�����xBƕ� (5I�!��Rn;�Ӯ-���d��=���ϐ�L)X�e�;TapGsI��0Վ�����T����q����,���XpY5��'(+��M,����ű1��ۼ�Y��)���M�֛���8�z*0��������Ɏ?��yg]�ά\l�a��n8������1Z�.��^I��hH�����k��~}�4�LUS#?�k$e
���ԦnkfÔ�7E��v->����v����%2�Lg�akAR��Ժ�T�>�١E�V��%`�rp?����V�m���6���:����!��$*�8�Λ4�I�ׯ]{��ve�tP{7����x�,)`�=x��3<O���br��ٽۛ�b�����$�OK���^ǪR���J��&[�Y>����/���sۏG-����2�Ԫ6���ݻ���뤑�����uF�UQ2{r���a���j,��ڻ唜 ���p�����B3!f�9��*�1�&ވElPx�g�C��!�Y��ky����`��G���=?�v���]R�E������%�"�5����	��X�9�_?u�j7�}��N�c��ΝdY���
$@��,w�Ճ3�+)]�Ϛ8�c��JD�{xy}�H����U�`4�Ņ� �
�]��J9����8v�q�B>�,��ǧP�����+�jX��!���[T������Ք�p��lb�������_��t����o2���:)��u��Iy��M�9r�}N�ƾ}7� �`���Ħ���vS�ś
��Ê�^2����e�}#0`?�	-Yw��l���b�	�����qӂ�+V�����ij�g|
a�ku�H`�	D�v`%;?=��|3O���8p�4)|��1����<p��X{��1Xw6ɩ�).Hp�{�_�)s�ia��e~0�=F��7l��������<�PX�w���(�����v\z,��Z������I�-_b��������
0�& %����&���nb�������T�yu���wOٳ!{�n>|��@�R��^�S�վ�<`�.�(�e��K�����pϝk
���~�����Zປ�`�yk��~�)�St��נ_U=4���yq���m�c���<��k�V�t���Q�k��g4�U�|���AO�Ӟ�y�x�qb�~ٓE9�S���:4�M�Ǹ���v~�ߍBv��@��vf񖋍}��[�W�_,�/ZP+Ѳ�,Ӗ���C�mOSR*i$�ŃC.���E��'!!��W�Wg�m�� �h��U�pO���{\�/�e���JM�8�W%&\Y������=�� %HpE�W� ���{��e+V���!��`�>X=���<>
&O�\Ѯ8���<f��5�t�4�7�����=m����5��#!xVT����>5�C4I����:��(�8s����4�9�o�:��1����}]�(�G<1+�ēZ�l��<Wѧ��8<��=y<���hj:����s?����%o�b4N��W���@t*���s��*�����6Rn��F��V}{q�'������Ϗ����*��&�|���Zk���AhZ�ʹҠd��yQQ�(К��� �]B*�:�}B$�-_�.{H!P��4���h�B����o��}�8�����5 �����U&3ж�ݻwx��5L`��E�Y���.:X���f�!F��4Ԧ��w����]����n7n��C�HUbJPY�N�~����B�?�&�Ǔ 2�����/�TM?q=l���c2��G���AK�pdz�|#���F�)���g!��H�E�
�繀�td	�����|<mz3tKߩe�L%c�JU����N.ʶ����S�<bbҜ�c�	HӼ� �� �n�{?kS�ǐ��ϟ�1��_�Ǔ 0x���ؿy��[�zO+���'�c � (]�>Q-k�435��؍��0�R]���� 7B� ���>~TG��K9 ��68�o��'^u�%?Ȯ(<U�-��7�v�T��A��6�(��n9�h�4��x��~x�`W�kqSq�>==�PҖa�"Q�����`����(����t~�"�	i�z~�,g�еrG,*8�K:��5/]���d r;4�=�yu�r���č-�[��wf9�7�(���Ѓ�K���yR{/�H�3�y�rk55�of}>�����W�����x��\�`�����}��~�i��j��S���|��e>�gKU�~���-�LY�z\\�
�������x{£����Z�����}8H;J�֡Px�yv����L������� �P�t�8��l0e����3���b�UT>�w~��Fa���QP��,xZS`f`��d<�ϾE�hM��"Ţ�.�?�fR+��6�n��6i�&�Ƃx�`طo�ቹ�����T���T�˜`{��h���Ϟ��fi{yz~ĳ] ���������K>�����pܤ���w�ǟ6��y;��k[��B�f.W��p�I+�����Z����1���z�5��!"��;��osj����IŤg7e�A���ԕ���?��bt kh��%�nb�9AK(�Q�M�?�>��<8��@k����OE�G� 8�]���=�f7��eSxT�S�������6δ����{ŪU� bn\����K�݁Pi0���V$% �M�k�:Y�։��מ}ef���U�}[��w���z��=`��bYكQ�� ��ͶZx����?���ǩ	�¢�՚K��9���;�]���~˾�F�oPN��~�?�Hv�*��_3�Օk���qK�/?V�������������[���ܼ�G�A��@!0h+��YV����-_�bÆ/����o�PU�����f�h�t ���_��v��g�dL��i��+��q�O���K��� ;��4MJ�u(��n�Y3o����w5�v��nB~ۚа���*~���q�ʹ�r(�'N�;�d�n���2���U�u��?�q�	���:pnM	�b�֊/2��DF��ч �K�NY��47���kj�x愞�`��\��?��zzy�0�|R���&@�;�[�qo�S�N
R���7�6^AM���D�>G�W �6@��a���B�խI����>$��t�=��խ:·���a��N�s�`��X���q��u�'�O����h�Y�d��Y�k���jyH�uʬ������Z��v�)|%�p����W� 5�-����v3f��� �o
��˱���ׯ�z��+�F<.�	n�Y�\),,�����|��EeǎBHSş?��d�xw]�$>uu������q��Nĩ�d]]K�U���/m��z׵{�*�]D&i�������a�4��u�~�m�b.͔�
���CL���U��|WAD|%S�\��Vj_�����4>������]����x<�.qme��x�~�9�@��f����.�2v�l)舘�?+���������pφq��<��"&oL�1Sӂ?]ͧ��"nϵAdC
&����Z�^ԋ6�z�o�>v�g� ���1ه$j	6�$�z��Œ�Z}q0Ѽ:c���N� �|�ڋ�眚��n/c��,ËǬ:�L�h��ڵkM�&ڑ5Yj��`1��22�! ��j໔��?0���8Z_��#4
�Ԑ��Ԏ�.�#iW��­�S3&ؗPyY�N>�k�z�"���;wV�������߉7���l[D�Z�߂X��l!���X�y��825W�I�����3_��0X9e���w��p������|�Gr:�m۶jp��ddF�',_{SL'�D@I�^�:{6��C�>]P�*�e�\��P�����rmc���Q�O hB{��@��S�ܞ
��yb�X�m�=���,D��ip.�퐬�؆��死�����A��vߗ;�:o��[TG� �
�n�t��g�� ���eq�Xى���e����Z��S��r�.T��`p��=��S[wם�={���P�hkC�c�b�˩�����6������� #�
l���	�b�D�)�����5��h:�q�<�W�XDH�̤^>p�T-v����`�5��������[g�a~���f�<�hձ:7�����a0+�-ˀ'(�������z����~Ygdeu*-!�)LC��U���'�V��wv���������bbb;f��;^����:?� ��c�܉�f����W��*��y?��u�R���h��SڙqL&��v�����c��¥o^�L�'U]˙�W9g$�E�����B0 ҙ5��rL�.
�����c����G��Ύ�s�}ʔ)��"��KCv t�ߟ��������V��ާ��$a���D����ѩ����H|'3����p2�P���b���u�?y"�{[b��(,��h� �x5��2��B��`*@�Hg�?�=~�ȩ-9t_�V�˗%��Fgݸv�F�G���3/�q��Sܬ�k�eP#~�����׹x��U0;��B�^�x�e��{u����d���r��#G c�A3��@D�:w�V�w�`8����cvc&��W:��OY�y6O�����Um�2%q�$�;�\RƟ@�w9�_���V���l>����|�!���9�]gv�fY�)����9\�"A���s欳oե;¸J6�MD6�-��y%�:1n��HK>:��Kٻ]�VrW����Æ����y����f�$���7:�L��a�,�����pr�huW���J(��j�yaЗ�l���E�?����f]0d��ӧ��%E��(�!�k��ǳc��O�=UQ����yx@�Џʽ���+��@�d_P���G��s�n�Ԛ���7(z�p�����. 3CJ��%�g����}{���GD��߿+i��P�׽��,G�}�a2�%�h\ !!�g�͞=�jҠ\i��W����K6L6�������<��!a9s7n[�S�S�E�0τӅ֧O�_R�;w���WSy|ܜ�qĳg�@��s��s��ޡD>x]j�P�����VS5���4�ҷX���E�	�ׇ���mgd+FF��[�n#���iXtW�%M�4��V�y�`�o=�s_&,l�Jn9~����[� ��8�p͉�ǎ=Er����XiޠnT-�x�
�mZ���U��(�q��\?߭���mU�fF��z�S�1�UϿ�R��,d�_����';�׹	�'?�Ȅ�ޓjGiظB79n�l[H�o]���o�6ڮ��tz0��#Ȉ[-c������ �}��S��g�c1sw���?���.#m���[��C�n�}��|T���i_�fBrg�,��H��ܢo�Q��H�ٵ�r�y��`[W���~?n�34�'��6��1�x�����+V<��5z8��m��S�a<Y��������i�i�[�I������e�9�x���KS���!�0�!c~���n��K9�_;T����V$+_�_�s�}6l�+:ѱ���i6�t�T �Ӽ\�sn��Ea��Q�D���3�&	:͔�u�u�V��+��ʝz�6�z��j��Ӹu�Lj��9%#�k\o|g,Nv�n����{n7C�RV]����@��>??t�42 ��
�V�e{z����#@>��	ʖ�df*1"_��*��g�0�kO�܏����;�r ß���?��a^BBB�|�����%9����-�2P@O��Iگ�����P��3�ڽoz;�������*<}�w$t��3�K6���t���w�
���:�b��ԉ�552Qlt�ه�m�	��18͕�yc,M<ΝO��ē-��,�dY!b�FYC>0_7D5nܿ�vhS�
`��܅��ƒ����Ɲ;a��G��ߓ��Ϝqr`�u�`'�|�dS �8����޿Wi^:0�� �qE�$��	`wEס����ܪEBB�1�ut�2�/k����D[�&g礋�<�)�q����`���/bsp[�ɖ�<�6&_�:V��C`j�ګ_�A�@��]�q�%9��:�G�/����U �י�-y�I��	�?��c���,n'�'�9�������ۘq�:�|{���^�39�?��J�7=�ڠ@O{�]��U���2��ω��y��o+�sf�;��_�&3�����L*BeK�ʁ3���;ʒ��q�`�N�b���ڎ���EnD`&Y�������/����] 5�#�w��Q���$ӟ�?�ό����o�����d�g�꽺%��L��۷$��;g��C5�^e��8�a�IC$m[+  ����V����X���a��~dc������zKXN*��0�k0X���Z!&���5���*.�3n����={����ot�
׎�`��S-�t[�I�-R�&9P�� 
h֓���M�����&Qp9HHH��A�BBC%c'�A7�c����S��E���w755��nT���IЗ_�p���u�	6&��0�0�ɐ3CSΘ1k�	Mf��t����?���y�r�����m��D����J_�\�	F��D�'����}vkӊ�B���QWI �ǆI�<=��+��b*�˲��y `���j�u�%���Ar�4�!=v���';ٱK��6�N`�V��xVS�̺{<������w��*�
$��L�i��-�� >PE�ӱ��)���H�'U/ ��S��%�E�A�?��M�_bL��z:�ß>U��� �ǞQ�wr���
��@MУ��A_d�2 �bgψ}���L�ԯG��A.��j�7hpFWɚ�#�{:p(��)?@6�h߾}aЖv���O��m��22N��w��kZ�_�X�u� �'�[�0��#��E#��ה����ȡ�S<}�b���x~;�q�ȸ��k�u�D�.����-��S�Q��۶�k���`H�$��+fj�@hK�Qw�ĵ$�,�͛ϒW�HPTE	/[&**�cܤ��GE�:ވ|�B��ix�8>�e;��)����Ԯ������O�Xr?�����VWE�z{�'�evF�[�?_*(�����*n���f������:�^�lY��}�����X�S[k�������1p����sA4���Z�T4�t7/36#ooo����T�nk�`�.��Yfܦ�g���ysi�p,H�f�}E���pd����&E�{���<:��U@��������g��ЅV+j�ί[;6���p�d������pP5�G�$��^Ob:�.�ɮ[1������2'�D����-	�8g�(JZe����o.���p�N�4|ch�L�X�;ͬ�]�VY~  ��|��Wu��CB+�v�tYҩR�fN���js���&�&Ӯg���}t6�_1�<�O�ۧ�1�6����������*O�荤��BxS=��ÿ�E��-��3p�T}߾��]HM<��}�0����%�7�Ywu������ݤ�̴��b�#��MǑ	�Z�$�� �w;��l���}{8koJ"�"8ʘ{roc�/ٲ�9.Y
���:4Р`��6m3���+��6��}՗Ⱥ�J���k�욅�Ϛ?�cz`X���M^Êk�Zq^:��;�����������惍~���YSE��ʗ�ы��"�_�Y�Q�|/�%�z?�q��js;��2_�!���w�[<+m~un!v%6`,��+�d�ee�w�����tNPj��e���Y����#���{����K����͈�����m���}�/(8\�sr^ ΐy�~Ta�h�A�j��>۾M�$q�v�!?�֯Yi�,��s��:���˗��"g�^�z;  ���j>w��a��b9/��;w�8U�x�����0��������R�Y:P2:�;���>>�
?�\�SWW7�����\o���%����w��a�b�fYYY����
��ۆ�=�������\K]����b
J�7o���-�%�%�Wz�+k2�tt��`dLptr2���`.^�u��x�|�[###��0D�D<�R�4���5�Ӭ�j��8��{v_�U`�ƍ_гm��D�Ca���D;b�v��:`��kɼ6n>x�U]��O�Cg�Y��=Ĵ#�++�����;:�,_��u�^�o��9��GEI�k��B��J�Y��J��O�x�#����������I�����k��f�9-���}]Y���zd.l>_��V�$wW[|��� RH]GQ[lV]Q��$��iR�4ntJ�}ک�8� i���N��	����h�8�U�"��x��߻{z�js��x�ζ��4"��#�||7�X7�yÌ�3cH���γI�����4-,,�EDA{��}�������yL�ͥ,c;�u'M"?Vǭ����)ph������?->��W���Q����A�:��"xՃ�?*���C/q�Z/%ţ������8����{_�p�������yy��s~�����˭ ��%a�M�QMSo�S`X�UQ�h�n���*,�~}����:�$�ȉ�$���I��n��rr��������!//��H�t�?�HmSq8�����R/_�ZP��C�ccei9K;J����*R� 	��|||��T�\�
���Ne��ŋ��W����:9�� �D/q0���]Q>o%|*�EBţ�9:�� (��%�� ���q���9�D��/�� ������>��d�n3=%Fuo&���H��(�-��g0�V��Z��(�X �@\�,����>3�:��+��y��R�Ι3'�;��B!��h�=��93�����&�GY�bHm��Mu�H]V�`[-a2"	�����>��g��m�ܮLnޭ��	̋�h{�`��m��tV�I|�2۾�����^\|�q~bUA���O���� �jAp.� ��ݸ�"�^}�*����2N7���a$	6��G�8���(�plq+��{��C�c2����{ g�����UA�NHH ?�xc����rBQ���l`}���kj�S�NÞ�Z�w��ԣsN�M'�i���Gl��ԉ
�cqw��D��\/�2�'���nՐ���%���[+RNˮ��Bۯ��\��g�2�! ���P8Afhݦ.G�0�5Z{+-�4H`0Y��sy�����%h���?��F&&tB���-��8a�4���w8���{O�Y�O~~{�U��b���$� ���CrsM�E��w�z��	��)}�!ɱkc�U�A���q��V�0�)��ymT
�>V��ս���ǌ��Q�;䬎ގ:�c�,�� �����ۃ=�IY(��%$&�^s��Ɩ��lG#l������!7����� 0-�%-����I�]{��w��8�ǧR��Ht��e'�&r��{�\��m.y�'O��u��ۜ�?.�D��ǲlŮ����J�V&S���������,Z�ڂ��=8 Q}#33ӐP�j]��\�M�N2+
1�T���mW)	�<AZ�	�MH�R���O�>1�֐	~�薟�ѡC�ɳ����"��D�w���:>��)[|l���s����#��@?��;鈱��L>y�ۼ�B�	���
�|a�����E?~���1��0�c�I��ӵ|�`L�`�B���_�~����`�#��w���ף��n�ُ���|����7����9�vJ�'�����1}YN��eA�z��F����sss�6n!�4Z�]tw�]�ќ�ZfB�������J
 ?��%TQGG�?&��15�R�2!cI��d��~�	AC��ׯ_z�1��C��	Љ�Pd���ݭ��$?���f@�*^ٯ&C5���>����٤���B)C�� �v�!CC.���d�kFOQ�Up ���M�{ɸq�P���	�\Y�G�Ⰴ4�'�:\S:��R�f%q��~,-��r�I�TK�4)����.2ȍw���`2���|�ʹ���R;4�?����cbb�Ga�
:%�Ç]�#��f����WD�Ir�+��`�� �2�������a$���NII�몡(���V��#�lqCcFz�Vf���r�����(|�h���"�`0�6��=�"��Q�� �0�L����Ю7Z�;wY>� �t��u�rG��J�Vx�g��H?�X���� �Ç�B�f�؃\�T&4���dd<_�~��F ��c�m#�d"w  ?WU�S����U�}9�c$޻9++��㔗e!���J-�l��D�'Yk,(!�8�|�כ<-4M����q&������87*z{ ;0}l#�a"�'�Me��oc%��֯V�@z��_�p!��!�oSKOKS������&���ǥN�V?��w��ڮ�;��ܷ#J��P@�k����� �*Ňw�𖖣|X�ה)8�+�]X[T^X�!���9����u�=�����2����� �'�8���3CHgq�uD����8�|�����J������?�s� 6�ڳ�����!���ק��+�e�Kd��h��;��3ٲ/_.�e�����Ə5g��y�ܐ���i���@���O@��8��o{2����p�<���6:Rwjֵ"e�1��_/,,���g���s�οr�VMk�7��$���
cAs�i���5`����tP�8{&�@�r2��6.�|N�;��lll�SS)�[����9Bly������

ϛa��/y���ђ����
i ����Z�.$�ʺ��k�8��I/�l�I���l�+-o#�Ɇ'��%��&�HD~������0�>ʾ�b�Q��',#OH���M�p�:�d�AS����,=�����{��Af �F�ۼ�\?`�i����y�7lB�8�T����x9�#���Y!!!������7H6����I�,�Z#��6� �U�d��dr��Y�4�� �?�]t,�y�:Y��&Mb�x:Zl6<���l-��Gx�����RR��<<OlĆ7��+.����S)��a���5�!��8����
]�d	��ȒO����x��>#�������~an'>d�X����G�j���]A�&\�aܞ@yo���4*�ʯ�����ܾ};��v������I
IzJ��Ya$Yo6s�ݨ6�^���N�.E��^t�׼�W�nS��er?@���{mIx�z�?����pa� �tǪ�z�! ۦN�J{f~��rcU�uw�����J�}�"%E�����;��,��}Y�e	2.[ir7�/t{�BdE6��lsu-����@O �О���m��*G��/(���k�US`���xPVZڃ�ܬ�-�
�};LnQTf��?����ܝV/�-]/���7�T6vj<0·_���l/߿��Xyl���~����Ĵ�M=p�!?0�٤�2�Lˇ�e�7H���:�;}����P���� ��@�G؛_ ��8���͕���1	ڴ�KRR�z2P�H6�a$]�����>���@�M����y�4��4��ܿ�|�N	�<@�]Փ>|�p�D!j2�����䙓\��T5���!����utXQ��� τ��X|=Z�}#"0�,*��a��Y8)��!�nޤl�M����dnvb�n�ȭ�����Q���^}�Օxp����ow�J\��F�L<�S���F��^ǿ�u}��^s���c9C?Ɂ!\�Rhʡ��O	\d1�}�����i�>Mz�Y�C�dD�8��6���p"�����<��f�KL�S#�^�%ƄA�3K�x_z`T��v�J(���<h:�yk:b#q<m:}��`������c�^�b& ��aDq%�[XD��X7�q�&c����d�|ڙFk�QQ;��9:)ɟLk��e�9���Ҷq��#��z�@b�:*GYK1!'��s_��>E�8h'F�^����V��';r����dtW<�N�~E�m��"/	�7#�^�,��|n�Hi�y+�N�Y Q&�r�jڇ+8��ۗ���2"�X��*�����nb��`z䱇�cy�9��5�c��a���|��R5�zY� w�$%-�\��XS�%�O�":�(�e�,�Yz!"Sȉ�n3l--g͙3��P/�v�{����6-���^j>�dl"Ȇ_@ ���2b�w��i���
2S�|��G�)m������C�e�-�#G���5�ó0up�L�FD�X+�$\I���IL�ވ�y�æ�"� HI�!�5��VP��0�^����l÷o�R7W|Gzuz%K��/>6�
ÊE��q�YRf�(���`&J��a~�xzMSr0A�8"�
�	�8{O �A>�����A-"���իL�N@��c qV��xq�t��D�St�Ӽ��Ԋ*գ!F�����::"���w�K[@���F�PP�50?�H��{���k��AJ1NuC/$��H�6���A�06C@U1C�D�ā�dw���.�g~o ���\����`��aMŸ������Y	���o:�'��CbT|�?�Z��DB����\K��ҽH�q�Q��[�⧹õ�W�C:e�b$̓�����1A���Yd�1u'%`tsĘ���ط���pYZ������4y��7��4AlS�Pr�'h����/�!!+U���[[Op�k��r���@'����@�v��h�'�ȓKJJ(rn�7�2�O�������ØF��yvgC>���*d�p��/m����J�N�3�M;|���0�Yd)��i;��4u��j�Oa�B��P����t`F?[[��������`Y%%�t���͵p��#��[�:��Ӟ�7�2�p�I�f~!~�T��>u��ڙ
�d�v!��P0�r��U��t0��'�h,�/���kuJ�_8P6�P�O��[zZ��?~��K��S��^�k��Wm,,M���3�{�0WYYY�;�W'���ꒃ�� ����T��၆�?)���?��ZǍg�I�������Xv�f��X�.H�_�g0�u��UPХ��ց>�~�@oCn���$<=�
�K�]������	�llk�8D����@�~�|���:�+t*&�%�T:u��'�:�\�����3�	�X9�z'��T��`�6c!B�d��H����܌��!��r��M���$���>��� �t8�ӝ�|�1����:���':[��WV�#L�+C�TЁ���k	�*4�j����spx?����0$-$���w����m��}ȍd������ ��G�o)�_sG����V����R<�N��jhjm��WA���TҬ��P�$�LJjĳR�s1����mUC-U�����<��jӭ����B������k�o� �UC�]�r�;�t��v�ܺ5��[ɍ647�����C�tmTT���*�@wKGw.��ܷ�|y/_�?"��U.��1���*��燿zp4:x������o��������;�-�ijqmR?����1�.����y�fB�+>#���zw-��"r���A�ܠ����5���~/�	�ZJ���yc���WG���ѩx���$�#SW\ƣ�x�D�:8�E�+��R�\��|��ׯ�iN��C,q'��#�nxx�mT��xx�BH�&+Vi������Ye�tp)Dd��[�����6���4�[��ꌝŪ���2(cGP$0L=lk���z���T\�L|�j�Pm���.]B�����^R?+� �S��%���}�H[;???��/�Z!23rdf@�]�!��Gs强�`�Տ��P��� 0Ćh�sCR#��w{��ؔ��{��[��*����X�j�$�>�ű�n9��Lw�^	gg�Jw��ɜ����	�|����2��]==Yqf�BB��&���I_c��0}�$�Uv��O�M����&-.��*�T�r:m�a��������u��h(�@�?�Vd}Uי����� )��9q�Whɒ%\\�lv#���y6/��o�����+s�C���4��<<< 83�>��.?���p��!tSP��2rv��r���$0����%����"�I�Cz��=Yi!/��������wSeP�*!E������p;�2�j�T�R��(�δ��E��N�/:�q�С��}4��g_FF�&2ϫ��0�lh��h ;)�g�Q�̾��+
6/N�o}�vtl�!i��~��.冑�T�A�T�wO�B�$��3+s����^�5Y��H�v i`�Jx��k��E&�U���Ν��˅)�;�������SQś�YT�x�+"L�O'��q8+Ng�ŋg�����̎���y�T��\���gd!�����$q���#�n�H�SRV�S���̝��%C����� �Bɴ.�#��{�����|*.�6p�ۺu 3Q2���4�H1jg�ND&����G<����Ɇ��g�k3�b?Lq�YBjtF��͜�'�� � T��F�/N�{������q��z����<����J�@_'u��nb��cqf��2�51<%���+8S�� �c�z'''�4V���`���Wm�!L���=�,�Cf�����T	i��Ǒ֗�b%P��L�pCxp����,[�SS��S���+�
����J���� �@u��߸�~���� H�H����=���H�	�gf���3gΐ��@���Ơ4:���P6;�H�����3�H<����`dD.���Lx�9���n��˾������ޒ'�+:��޻}����Y�w����)n���`ߊ�OJ��V܄�G��a�)^��y���ԃ�++UITZ>���!-_)��ިǡ��C=����^N}mj�����ʾ_���{�ʑ/�b�
��5���M�FL$OL���R^D�<��g
fv5�j�� [D�����tk<���˒>}��(�sqU,{� �Rq��q:��I����,���i?pqϤ�c?�J�W4`v
~ͬ����'O��yYn��S)����ԶR�Z�.Xx��̊1ɗ�$Y��b�`^�쥥#n���]k�bɠ> czSӱiӦm/�����\V�i��yai)υ��$EyYW�r�%���Չ"ҝa�[� ��އH�����j������|�J+W�L�[e���
���f�����W�
�e�$�[���?�g���m���	����b������RDĪ�t��n�%�gY[��K�R,�\�U��������P΋��ڡ��'O�~�1��������s�H{��^@�S[�G@"������@���,4]khg���s�^ �ܝ��V����xh:�
�B��D��9�0z>.�����S*��+xxx�����e����r��ܹS��A�ғ�<$����v�Y\����?�����M72������2H�1�9��v���n$Ҥ������3�=mʷ�D?޾��7V�:j�4{Bj����� � l�"��1]���i��}��u�;��8_����v}��8�=��IHH��F?�1���贡4�����
�DGGs�t -���J�����SwO�](��@��@ ����W`՗/_;�b��冠Du"J�\�lJ�aLF�/\�_�-F,/��#�����ۊ��á�m��%w��Rnr&�L��%|�(�IB^^���xײM���΃]�V���e>��s qPpY�����q�C�ya�CKKK���dH���TBԛ�ʿno��땱_G������.X�KJZ�$ws�yg�q�C�E��%�`k{�������Fx�n�������k�_/w���7�ȄA%k�H��V�E�T�eJ`�/L�w�q��	��э��<���va����K2�ow�����Q{E�ߺϬ#ٮw,�%qi����0jp�u�544p'�3����6��T�90������\�hϕ��
3pM�u�(3.L�]���^�߀�(�ejj !���G(��2~~~��k�&͛7O�ak��-D䤧o=~�Rx�
���J[��[X���o*Z^<(���1��z���V�p	��,�.�- okK���S����Ex���D����Cbbb�l�r��'��!�}ŎJk�QN<�p�^��g/K���
�|�n7ߗ;5�������A ���ń�^i�z��5�[�������m��H�Ǐ�.HP
�hB���$ˋ�ES����f��������J���$�֊K����_��'Ӱ�_@ ��ʹH맺�7�㥑�	�9���9�7�Ν���#{��g&��ų���NЛM��ᅦ�{o<*Oi ���~����NL�+�p}-����@��=��߿?~@8F .Cf�"���+�N�UV²���~��-.�{����{K�Y`Hc�Θ�-��~j��H�_?����a�M���Y��50����&����#3��}!��M����ԩ�g�1�)*,,̡�ۜ�ǲ������B2����|�J#A�B��]��7߿���`�c��ϭBFZ�*���=qCg3w��y���#��k�B|�"���KjjQ�ی&pW$qgpee����{�� �ҷ�6�ޓ�����K>�����y�H\
}�oG�'��m�2�����+�ŗGn8h]RZZ�Vg��0#'�mϾ��{��x�(�~*�	�n}�n(a7�Չ@�r�B0������!e��ޣ{s��x���/_�z����;� �­��
>]]]H.HG�c=�}��/+�
���Ms�ҙ<b����/y�U��^t�������j�;K�+����Az�����vS̿���Tأk�R���#)))!)9b�Rt��c��۷�����>�?��.2�r+n��Ua�����X\��WÞ#�7- >9�O� ����z))�
nS�ٗ*��~H{��(BE^�S�G����ց_�Z@�^��h��^GSq��@�ճg϶�|�E��8��J�)x"3�
��Z�d������U�~Y�Wi��nݺU��S(�}^pjY\��^Fx���� �Y&�{x�Q��o�����Ǐ��˙I�A�m��Ȕj�'$[�����/y��	��вEO��A^�����B���e%���W��S<(22��OsTU����)p����@""�`r=��9�����%ɵ����;�{���JԞ.�2Vj) 5p�[w�I���0�v���ڸ����̮銅����=�a~o�%.C}�2��?L �@�{��h�h�c�����4==.V@�/y�231F�<��H��I��{<���ɠ�__��^���6]���n�$*
��xP��8��Ç��I�&����̕������J��0�9tq���ԝhSAjF�`L��P���� ��^PP�_�u H�緵��Lܥ	9#�z��yվ�G��遌�}]M��hj҉����cK�����~�b6d�B�
����3�����$�X�OP�}O��6�z
���Gu������%������ҫ1��ON��^�0<�y����`E`9H�K�&�U��ؑ��@�Ģ�QI�:���6��e}�n��a�˸8n��	Q�A|:q�������?�������Pd���S���C<4�ĔQf<Ŕ<!9�LpѦ��d��W�����/".*�D���8���\ӂ}X;��{�3�&���p���|�Q �dn�
(O�;)P�]!�Pi���Z��_{HII)m�{��?��[l.��3Oo%D���ϧO�p�6�CR[c�(��իW	*�4'9�������� q2?��1:z���A����߈?qqq|0M�/_��a'�Q���jA�H��,�7�#�׻BԪ���g�<9{�%���:�lmo�>Ev�m�i��ў�{\P��b-"��u<U��,f��+L�տd����E!t[����؅�T؟v�a>{��3D���� �%д���{�@�[���:�o}�jFvvv�����uƠ������O󉉉�'/�:�%��TC�l�Mzn�/-�ꪭ5V%�2Q|_����-T�����{�D'�-�X9����^���!�X�����3w����/C$%�d㬥��=6/�ͭ�2��.|��D�c�+�ou�����O���!�~С� �'�$,�_����ܼ3`�I�[�V*��ٍ�eUU��޽jd�H6��.@3��߈��D�D(��)ݹsg$[8�>D):
��N��_�� W�6sfh���$��
__ߺ�p�K^�����l>���"��a��C��W=�ƍ��d���Ӯ-�8�f�����L�V87�H�����ee*$O^�'z�l�c�I(͵��?I��R�UVN��͛7ӷm%o>'յ��ߘ#�&UH�ه�`�n�����U)�C]�����os�^Gin�y ����1��+8�=Eu�ɠ|ҷ97�5ku��Y��R���QytQ�H6��ս�~�GUg�R� BK��R��%6���+c���/��\Y ȩ�r������R+���Ç鵵ɡ�i!�m�f�J��(U�?~���.��������G*�g�! 䅟�no�9�]�x��m髵+JKK��t���
\h`���!ₚ"��!��laH��7-��d���挌���a��~�J&M�D_5�~>X��|��M-MӲ�-R���J��^�!�A��򆆆BZZZ��]P�$��aWK�Y3+888L2h�-'�F��}�cx���U�.6ia$�������w�;wwg��4s����,'߾������!�#t W /ڦ�&��tCȗW�e?��X������O^9��Z���� `�����[��A^� ���(�*SA������}w�S�84��`y��kn�E����F�d��RqƊ6�]+#ww���|�,@0 �I�n�_	���Qh�X����	z�K)�*�#���$�È��}F�t���̭�y�^���u�	��9o��	I�Uǭv `GfM�sT�ޑ���QQ���@�_��aem}������1K��.@1F|e������e���C��`�g����kcq�'� B��w�(R����d�� F�݂�j�T5�=���jT�\�?���v��kJ��?c{|rK^dܸ�f��Յԇ)��a�K(�E��e��%P�뒙�T\颵c�nϨ�����c�A����wt����� 	�ydmou���k�i>ԏr2f5��:0h.��m�xE� + �qۙG:l��s��4ʵtU�Biǟ�fӵ|x/D�h˺���w����_��a�����gv�S����XB��?��X�_��٣n�y��]n�@���.��f�fy�����כ�<U_#d),8x	�pW��:ҁ_����[$���I�\�B�/_ޒq������YWl�q�V2�+ �q����|��1�bC:��nJC#d`c��@�	K��M1$&�.5^��[SSSě�
���JWrr ���(���� �e�T�%��N��+窞Y�� �����Hti;(�۷o{����6��|\�1��M����A �*�H���v�H;R������wV����+�H?� ��"R�C�3�4��U�͔���ѕ����,�w�������P��s94�S�H�/(.���b��iN�Gwh�s���������J��ʉ���{��ۂ���즴��uSR
���go9�n\�֠sHj;	XF�N�i�MMM�Q�C2XP�2�/�� F�"�B����G�/�Q�`w9M�θ��N
��?�
�窪=��X	2yD��y�R���&E1A�R.�jd_4��LI9����|��ގ/��M���_c�4�ƺF��-(��5�7I�F��ݳB��V&/��F����.������i�d�ñ�Dҭ���+���R�"U�<�� �W��m`�=�z�6t�RB�/wh��p��%�J�֑07�`̠e�qk��" $�TUq�>���O��I�աA�E��[n^��A�Y5̌���Q�n;��mĴ#i�5e������oR٨�vS%���sp���,�!D�v��m��o�����c��Jw/�dp/�7�(F.�`d)����>���u�Lʼ��S.l.:�N��O��� �����P�s��W��o����G�c��ڃR�嶗W	/�^�UJrfd;Y|3#��h^���{&y<4	��z��#�?z0����� `�Lo�;|x)��-3n{#~�0kS�;9�.���^D��v�6i�p.��'��$���ᮕ9/ȼFF>V}��p�B�,�&zQ�f$�
�$^�4��{��c��jL��OE�ѐQHE�
�}�eiA(K*�ڛk�Lbh!i�&٢�%4*KB�QR�M�^��s?�����ǌwzz������Z�йlC+���̷s�k����р#�[�;2�}�����W�-CD��رc�O�c?�
���S=��Ӥw��A^%�TU����0t|��F��nc��rF��N�p;OǕ
�i�ǔ������%�~�����#�L���zڞB��?��	%wH\�� b�����Oԗ=���*sbo��4u��o��UE���F���܏��q?*��l�q@�Y��dC]Kj�!�`.��lJ3A5#�^�*+A�u�z�j}i�~�����m��D�������āU8H�ߜw��\0 C��������k����l<:'f��3ڢ�he/�����☯<����AO0M��A��h me����r��pFMN��| O'�d]\�6�y������0��L��/0��鞿2�j�ѯ���2�1� <9>�T�V?G\sϞ=W�3`�d&�'!eEY�Tx1U�C�^Kr����P0ǝ����Y%n\�D'Ԑ�(~�?�}�_�,N�@�4E����9w���������A[�����%~�/�X 7��?������%԰8���q�)'�-�j����Y�*�On ���ܺc����/�V�>}��{i&�eecI�؀�Ay71��;�I� � b�dݮ���&�]G�����ի�|�hH�ќ�DXɕ�%a���"�^e"<y���yZ|�!ã�*X�����P>y��9c8���f��h��abO���jjj�����qz��c��K�C�����;w8�Ī
�"G7Q���~)ս�Aww�C� r��nO�Lqs����K����������)W�I�1a�����0�|���ZR�߄1F��ӧ�.5k��Y��0�ix�V�v�к	�5�	CW����U=�� ي�ݤ�t������ZڻW��ݒ���~����?Ҷ��&3�k~N��~xSmt�%�ձkq;��:�Κ5���z��6��(��������ܒ�ēGT�cB扃�����w��. j�Z������|C�N�uX"pK=����xWcf0�
}v#��̴�޷�fq���V��8����qt�W�J�����i���U��::?&�`P��)��x3����?��=�!���V�����&:GbI���7N�Hv[��hW�%�����rh�%��RR�����*�-۾�X���!C|��l;l�;��|>_Bv7x�"!@��ݱc,W&�0�^�7LƷ�����
n���<Mb/�W͡�D�Eb�n���-�E\�K�`��/�Q)���Z=4�x��ss���!cU>��;Nf/P��n���s�1��$:�לdU�.��G^��ZՌ�\N	�S� X��k֙\�%(�eqX��}��K�ݰ�b���0*&��e���g�2��GW.�k��3tu���L}��N�߼��>�:<���U=}�}����=���z��G��?v_�<�_�Zn����G�u��l����Q������3���.r7Y"w����J���S=�s��o�D�U�f}�B�y����K�7��Po��[Zj!;� �[��}�f���-=[�9�\��)K�O#����ĤA��[m'T���?[o�C�Pn�?r�&C'�c�l���N���3�HJ�{��\
Z[ˍm���֫��6��~��1%r��>O�c���V��WW��s�ނ�����޲�!�Ky_��&����R��gΜ��ii�d������7G�'�v(y�
Z���<��N��4��N/T����t�mW�c�2��U#�)l޶�mb�|ϖ��!�C�a�jP���ʰSiC-�a؊01�+���ϙ3g��7�"�v��%�����{�>�w�S�C��O��30�];����3�#$a�7ֶ |u���;z��6�]p�+����������rw��C�=Z�zuN��P��N�:����gmd	%��HOt��Ev���������<� Z�^��D��O��"�s˶�Du:C�����gۢ��?}���N�>"�u0����`ѧ�/)gd���}���V��$�C�xF�yﻌ�wC��M�3��>��������.'����q#���v�W����_�~����8��~�/��0&�db�v�٣V����O����9�724�v��?d)���a���'ҿw�Ћ�LW��Wׁ��+s�Ml�$0h;q�CJ�v� ��.�!-�K1T��09j7Վ�?^7"^8#��=�#=z�Qo��w=ЀO�܁)��UUU�{��4���3��8��G�GbD~����!�K6m��5c������o��v�[Kv���Y�F9��-���-O����7�m�f�3��BS^��}�	s|:].���*i�;�UZ��U&AO��������O㴽y�x�ոp�����j=� |����Û����W�-�Bs���o��֎u{������Ƃ�яM3S�AV
��M�&GVD�����8���f8T����}�� ��!![�P���1N�0((�5{rC�,;��^:���$7~�Ā���w�&N�4��2��.\h9���K�5��݆t�D�3c�?�pBR~7ww&1�e����7�d��`�⷗>�7aP8���ޔ�#�3&6G�����c�h�U�R d��D:��CJ�}}ǚ�-V�y��g��W��I��e�r�֭�2��� v	�K�N�b�@rώ-���7�<8�����-�Gz�N��_
�BTg_
��r*�T�}�]q�He�mo��mfI�Ro�ʂD���Z�Wan��� 9��X�2>�<}��ļ�y�ŧ�R�x�����0������8=������d��Q�>FV�4F<H$�TA�iL�rn���z1�a�>�����C'��vs(!I����X�ZM̠���f�Y�e�1��tJi��Fo���4�'U^=ń�Sn\��*k`=����Q��v
'z�tF(|S�y6��f�5(S~�Ϝ�ߕX'��[S_r�2�xpũ�OI��n�@��覿�:�P@\2�.2Nn߀`{~���㉳��)�����Wqr�ǫ�$�ǬGd�R�pq��L���P�[�p�Õ�����^,<�ӿ�$����M�(X�n�+�O�y�����v;��A$&��LLLL���`��l�֓yr��jy[w옴d�2���2*��o�l�;L�Ǌ��� �u�ɞ!�ʊ1�&���C�<�	zyz����_��F�.�}}:�w-�����y�s��S�"��n�$��wp�S݋X2)����IH��o�F HZ��᥅j��7�=��M�VI6�(��_t���?G�����B�������`�,g`�
�#e���&��]�qFN~�����إHг��W�NNA�e�^f��襱���QD$�]�un�F��V�h�M�Y��R'�~}��}�.�	���_N����c.���h���a~�����H�0��i�l�*m�,<$�����h0hРX�7�H��^L����!O�-���k���s[uc�qLF���� TB�X�(���!� 9$K~�Nv�';::��#�p����e��d�4z����>/R)����C�o@3�4���dDi�v5\P��!��i�^H�},N 4���M�n��[f����ӕ@��ڣ~C�Q������a�xZ���T�8���
|1��^߲�u!��#����z2��N��J�f��~Ii�qb�_�8�;��!IꨋK`ި�
`����Z<�-�wO��y��tӔ�����5��U"
�$�p3�%��SNǍ�g@�y�0=���yt%�G��m��_����ه�Oo��ܩ�oUY������\�p!�b��ÜS��PuK����@���+�O	�0cR���|w.'BU��KE�o��ǏW�ͅZ�f��N��T�;�	�#N�h7	P��Uo��Wv�JRfW���o�-�=MQ������5�\xkBj0������t ��x����l&�u����r}���t�]K�L�V(�eb����5"�h��7}����ya�tt�f�֯��<�X_oA��QzӾqP�;g�Fy�P�a�W�#OK����!TG^�����66UQ}�}�I			�@o�����+��� iyh~ľjq^�Ι3g_��n�	����aJ�����;w�.���GXa�ފ�29��Ed���nG��a:7��<+f��P���l� �M��a#j�����ER}x�SE_ϓ�}���Ƈ~��]@8ݫ���%`��t(<���9�e{\.��U>�:�d��?6�idf�z��qI�ٸ�Nه���?2�E1[�ƒ3AP�I��3oa��S���%[��b��*�?r�Ѹ��-�[�P���yLė?�&����h��'�uu�*z.J�������K�������U��L�lmU��D:4ϧ�>�vk?{��C��v�wz��Y�v \6�e4��%���,R\&���{-7h�lT�����1I��[&�����lq�,z┐$<h� ��S��U����K���&K���2{_�����J�J���74UE��j��ܯ���JTR���6�G�Z�����yռ0t��+�{K���qwMKG[oo��'�oذ��r!�\������4�Ɉr�h�����Sf+��svv��7X��k�O���q�c+�Te�� �Wv� ��ʭ"�le�ߖ`3��D E���K]ѝIi�.���%�d��r2�m	�>]w���5�5�#�FB��ˇD�������<'�����x�<4���L�����w��,����:y\�/d�Z�d{B���Tᒝ�������x���tYZ���ԅ��~5u�$ۧ2�#�Vd��!�\Z^�a_�(SMK�����S�"���6'��K���4v?�'J,�G ���8��OC{���̩�OeV�����r@0a}J�}E��(��~UZ��3:�Sjdv�`Vr��4q�Y��Ԫ���j��jE��Щo51�x���.��F �.3��JW�b��>?�[P��@jj*�~�>��7��q��L?B��&s�>M�yc��о�Z4n�u���;i�Qߤqğ�Hc�A���_T�۝P�{w��?ca"Fpn��}�4P�N6P�����٨��|�TE��i!�m�Mz��6ʶU�q1���=����{��i�[Ӽ�e��߀����ʮYP�p�0��K򕽟s�88���ZT������C0�Y+q�N����cB&kF�O�����Q�yϒ8�XBL�M�x����9�!�[���0�k�jk��a �(���#"����o��b��H���B�:�{¦��Z����(ciz{_���h�GӍfrvA�me>T����)v
�gU�'�}iff����H�HG��T�TJ�~] �6�xiW.,����������%.,�" 'V�7U ��6��YQ��455���ﵵͥ˭,{�~�7���ӧO��S.������R�>,n�}�(]pѐ��32�eҽ�Z��a����c�O*�}�U�ۂ�|��r�0#l^n�b�"
b��?]���C�-9�/ͺ۫�Q��lQSv�����Iv�l��L�,\jQ�9w���ܿ���h�����G�p�|&�p�$�t�7m�F���)U�X�;i���
�7��c������a���'����z����o���>ܘ٧G�	��i>��|�݋'7(E�."*�L��a��z�p��<������Ǝz�zC����"���dYC��B=&��T��7�E�e��a��bGs.��R��-�������t>~��Jp��Z�oP˙�Z�ʏ�!+~qͷ�|E�<�Y�RK��{���3d�א.���3�%�>���)�O�����n���z���T]Ku��������x��K;���/��+a3�*:�_�F%4����ɓ�B恒9bB���Mb�����}0�O7�Dj{Kmeؽ�;g]�q��,��ٮ���K*z�+��s�.��A��`cck�Gֶ���-[��N.�;Y�5|��ѕ���I��iHl�Ç����?@���>��>m46��\dOW[ɘ�U8�FD\��6k����[�,t�@���/�2gm�)�&MJ��\F�U0n�a\o?�}�>�0i��/��Cy<����5��G�7�I�龂r4�J�e"9��1Id��[��6�����o8eU��q^������7n�`_�}���k�Bd F#[�b~�Q'��Y�a��cǎ���k\���y~"�����FE@��^�|H�j��v��,����qX�5K�0�HW]�m�JRMK�-�x"����n�\�8�J�B�(��Ԍ�T!&Y��/���vRf$���T:K5�7R$
���,� ��9�9SKFr7Y�vl�p�狐��W�"׋�l�MMkn���� �CF����^%(2!	��/�E:�eC�A�&���� ����A|ѩ�����h���kgͻ7�!"n�&�Y�1������3{Y��V�Y$'�D��r�$<..���G/&�_3����x�˖�R������c*�`���1��m����6Ɵ���?
����MO^J�����%l�wu��c膂b 9r�Z.��^Y\h�����l���o��xv;�YwC�ߢ�S__���~L��e����PB�m�0�Xt!�f͚�ġT!�z�X	[x�G L��	��F�%��%-ӳ��JOO��n����ƪWH�X7dxP {S����)O"���g|���4rsK�R���q����C_����8����G'�����wւ����<a,�����[7��t�q���yR�f�m��̤$���IE�|�}=�s$�-LS�AͰ�pxX~�yBNdݮ��}Nr�ZB^�	�թ�����R�_��r��!�VV��n.��,�?��� ٸ��l�����D_&��� �r��U��� ������xW�	�	֙�5�ၤ����_���z����Lr={f���}� zŲ5s��e۾�ԐY��d�Z�Ur����Q����� 9f�ZosԂ*���Woq��{1y�b�]gy�������9��8g�dcDE��*��n�$��':�����Ĉv�vM�aD	��i������hw�T��ۉ�����	�/3�,�XĶV��_�@i"���s�,�S�}F^���ׅ����$��k�.�̈́b"(MJ�n�s42fۆQh�1�44sQ�:T4t!82t�ؑ1IJA.m��������}�$Ǭ�ap��n�]��W��q�EI�E~����YI�oo��*8L�P����NN�(е��n
ϿOs�LY�#c������ݯ� ����"�����L^�5��An;3Mb��+�A��(��:t��D�钮e�������E��a�\Xs�\�F�i~}���� �8k��%��؁)�]��]}�j�o��z�yL�V7�d6�����COT�l�͸���8ƝǻJ�?#����Bo1�.vR��9]�׌~��鹰�/M�C��U�V�C����bUg�AV��r��mu�7�]��1�EHo?4�6�%�0�i���b��2�,n1�S��h[C,,
��E�����+�:�[� �eo�s��!��٢H��*�CyM�� �,D���I�߿�L,� ����'�{���]���ڛ.�Aɋ+��{�P�5��ʽ�j���	
zqW��W3��3ȣ[��YOo���W�#W��d����z��F�'y4o��?����T��J��CI����Qس�'Z���G��F���hy�û�&�����:F�n��lj���dg�v�����W��׾�����1E>~�ݭ[�V�2��薫s`���7��<�4' �	:����<���H��}#����SbN�ԏN1wC w5,�n8����-O����l�n�CX�#�x㸈��ξ[�{�i����#?����uuGKHH�:�� 2���(RB:�X-�@DC����l�
Az��qIK���(M�v���:	$�z��/���b���Չ��x�
�3�7��2r�O+
�=>�[� �	6<��M���^���s?�̳�l�Ά8<��6�k��Ѯ濹T�m�$�!� 9K���FE.w��n�Z���;QH7��_T�\]]������Vk��C�2A����Y{'̸
����������K���=o6�����3UY�fe��1�8͹�%�x��f��ˮ~_fp�����ȓ�/sen�٭���z�V�_]I2����#v�|Ì��E�ˣ��#5F����q���lT���5�6s����99�G�J#9�I�����@>{ 94��WV�c��y���M�!Y�z����9=�D�"�>�����h�	�;��J��`�6g~\v�$/��$_,�M'֍�uǉ������U�*d*s�q�e�y
=����e�Gs�q�y�S���ows.i�������@��کd�J|ӏh|��e� 6L�>wx{w��e^�DiGK����.��~��C�m�D�B/�?�vNμ���fn����t���[�#�� ���l+�h�����5��Qd�Q�x����:��!�fl_����;P�<V� ��|^v�"������(�\�w��!��I�$���wC3�V�*(Fb"`7b_x�EZ/s�$�U�6�|U����i���+	���:�B!'Rc�z�qa4���q����%�{�E�7D�3���a����E�Lt��zG5���rLR̯���6Z��H`��_���D���K�_�]�x$!��W���Ɏp<�˼ܗa�C�:[w~�"�톊<���"fϷ����lUE��VT`ؽF�{�""��eh�n`A�Y�aL�`7��x�
ԡ�x�FF����II=h� �ߧNQ�O���7V=F��x��Ӣ��	.zq��Nn߀z=&dz����v~���ȟ�^�"Vy��:UY��hq9GO��z�q[H>jS3������Q�A��5�u῱r�u�5Q��^p�u���gn>՟�t��+W������^ed��M��g�Z���HN<	��X�����&v��L�v���������"�Q�q�DE��b27�����
}+��+����'Uº,�Z����@O���|����7��w��2�� b����#������>+� xfE���n&��z��+�,��'���#�����Q��Z�:�[a��ݱZ�V¶�@�ۄH��uڡ�@������۷" �HӲשd�Ǩ^\� ���M@#]Z��-ۂ���yu�I�lJ�s��:#��ȒN��*Ku�qu��Ә���o5�P�ej;lxȊ�����n-�w�#�h7Ë,��nC��йL�G�f���]i�
ݨ-)���gu]�uKF��l{!o7�$s�d�z;
��qUA�>r�$�.�Z��[0��Bv��׿Q�iY��Va�}�]
<�L!`,'|_=��0H�e���B��1&*M\�.I�bba�V0�m>�G�B^^��ll��eY��?��@4��\����P�&_���4�Ν;�x�}p�Gr*���"��R{�����7�_�o2oƕ���6@��֖����f�e��=i����}�|2�ꡦ5�ф���*����~\��J��i��Rc����ݣo��gǾ}3ԭ��!Ղ����ij��ِyvNN�Q.j�t�[�q�Y���d,�� ��C�>~;0P�kc���%N��-&���|��s�j��@4��j'"�`�!����?�`�>�PO1�"�*PAjM{�zyX�+t�,�i�Q�[����V�����pv{s�_�2����R�(�F�q۰GUUU��T.&�vH�wYX��俭�,�||�Yex3��t R ]a�����X���ȫ݌DY��(⨤�J���h�!:��=�u�,<J�{�d��5��� ��h�$��n��\�4`����aF$�4���{8=u��t���˥����'5�i�1aH�%.%��SW��N�7�$�C=(ݻ�Y�CO̱#�0c�\E�h=��6@��K���������b٢n�WWq�XҰ���ݞ�.ڨ��-��*�aW���1RCÃ�.�>����T`oo�S��g}7Ͼ~u���O{A�a��G�ApB�P&B!%%B���)�\���|�fN*P��	��5��ja2�U��Om5��[���X���A�I�\�@RK��9�@���w�l$͎R�L��(��]u�F�(#�b((��S��Kcvr�8�)dT������W"��14�k�9/�nٗro�l�k��Jʪod"���?�n��iň�������U�F�2v7���GM�O<�tL�-�``�鋷��^�"##k*0�6mZ�Υ��f�og-}UQ��đ�����Hc�l�
�P�u�8X�yV�y�1L���t~�����	�F�>̀�'ad�?��cz���\T|�lV���c,r��������)D8X0���-��A���2�Uͼ���r2������i8�,R��k�KɕՀͳ�M0�劘�8[5x��Uz��q�����^b�H�8Ѝ37!��GR��#���_�B7�E)�^��J>L�iB~�>Cĵ��tǸT���w��'X��ir�΂3:9��ŭ���r
�Ua8���Ή��A�"/�8?����x�h��P$�v�o���'���o'㦀k�g�9`�\ ��?�z�H�6ڑ�?T ���f��i�!3�a~�[��׫Qh�'����	Y5�9�$��)"k�S8#�����bbfc��Me�;���lfL�5y����	�('���+yc��. ؈*t����e)�����a�i8�^�$���e������1�]�vJ�|ڱ�<c�a^&;"�^�<{;�YY�CS �k��"(@�X$9�?�Fdj$��1�@
+�����Ɉ��O%�t��4FT��8T�I��t����S�l����LLv���5�t�����$���.���̟����ZܲUe���i�y�q�	�\{��H265�'A��I#��%R��	;�o�u����ZD*���,���m!�1�Ѥ��t���#ze�s���4���Rfo��Zn��Ek�pQ8�da�__�,)������
��h�H
;bt��x�M�oy7�~��w"�*,�3(F�e�*Aj׏f���G�j�o�}$\M7��2alZ{�������	䤥��+W��o�]s�����%������E��g�<H �@��q�Ü�^L6?}�pm��ג��хX�d�[�Q5Md�D"	��g(�_�cm$�@'\��2����O�ZO	A.��h�Z���Q�߾�yl��H&r�?�M�p��$�>�C���(U��i�E���儂�cF�-3摒���a_���{.�ӳ>�������c�K�Gha��M������f#�*�Ė��Z��C�=ʨ� <���~���4�Ԑ�e�ά-^��Ŋ^��ID)���WXZnurzZ@w�g#�U�K�K���1�}^��lKE�t���͕��44�:];%��W�n�JQ��S�"�3�@��o�$nĈxiz��t�}�]h;5y���� `�ŀ���.���M�&dA��K{L�j��.#�@@����QI���k�>��0K?F�g�pl�����X�ӯ_�r�O9�֐���,�7��.�	
�Ҳ���^����=������?�|_���ؤ�+5��ȶ,�c�E�|��.l��o�C󰂅}����P�S���i�30㎸:@�b����cp{c�X���!3����Kgl��#�S|{R�Z��"����M�a�-[�c�	�u�KPBF�Wq~���6���3۾�-J��.�5���x�%������vb��6����f�dK������@K�ƙ]e��b��HS|�+�r������|�ޚ��jM<$���JI�f��[����R�ˎ��M���Nk����=�qp�\�J���`��A�r�Α�QU���r>ɬ_�[ ���e̱�Ň�߭�s5אD�)�0Lw$A�k6ⲯ�ˑ`��z�~N��D�%%%�[a�1qVv\������y0�3�o��
��B^�e�\Ǿ��,7���j��e��ٚ3g�k����l�)
4��%��lx�ҩ��f�F�c�R�V$d��I
s�!���k���/�.�}���p8dQ����T/�0A_wD+��4���@�h�1�j2Sut`uğ3BV�J��`�%3��a3]�T#C������%d_�`� ����3]_8�1�G)���M���N�`ޓ�����㘂�NL��d3΀�l#6����4O0BhYCΐy��=�>]�w�K��g�s��Q�J�`a�HG@��l��t���6+�zcȞ7�v5"j�5�&�z������СC��/�J�{4�R@�.c==�Ɉ=�_O��b�z~�w�~\��T��%dk����d4�[+�u�D;���S��� �����x�ǎ�j���O5N���"-�� v�k�'����81dc��,(i���l�I���EHd[A�k�9���R^�zVs���nV�0x_t�-��F�g��}t1�Hz��d��oa���\��z�ԩS�e�dt���9�K���-S#і�j���[��6>������N�Y?LQx����'s͔�E��!t0��]^���c��c��+Αh3�j̯�W�@������E�Q#�ӣ�b�{��G��J����IKS��"U��L27��S��
�����U�p��!�(��Y���5��e��Lh�dE�F6}+�J,��LoHfx �+�z�8����DZ��'&�^�ӊX�XY偤��)���Oቄ�Xt����,T��[+�r���rߵ������*�݃����ҫ��W���[B����;g�t!��'N�ؤb灏�	�~~!�g͜)}:�`[��.���b�]=�kZ���C�G�}F�=3��\D����u���ȯ
Ƣ�`@h�>���0�{��߉�����q��X-?f�ʰ���|>~d'u�����},��𹌣�DY�A(a��*�^�q9H��<�
��R��j"�О
��B����S�,�#��Z�p!�q�˗/�^'Qsh0����#R�1JJ�cf�]��q�衁RC�;IE�L_�7��3(�h��iJh^����٠��GJ�`����ҍ��z*q����f�i�����n�c1�F�C��]o��fԺ	sM�l�L�ᕡ�9¶Ջ� ---�O���ʭ,���#�O',�)�cX��בg���2����H���
B����s��M<0�D~j�UK�f'�<R㣚�ve&s�B$�s�Z;�K���ݻ�����xjǓE�
9M�aaA��=��r�ΝQ>_�-��L�`�n���F�
�E��mG�9|�XVk&��ӱ	�v�:������E�$2��Q<|�\!�����I`5n��t�)�cUk������t��8]�Z�"s����<�V����DW��\��2_����l��Tﵢ]ц**���Œǖ����(���YgT�?�"��FF�FByI���[��~S��s����^��Z�_a|��?����޴���6?�F�>L;���ܹuR�?rb�)*��X��#�CH&�a%K����B�I���&��#��Ѥ�X)�vJ�V����e�b2���Y�9�3k0\�ng��I�܂���`�wm��{��7��:j�˘�*�t���_ì�X����^6��q(V<��x���I[Ko��m��މ��Z�~�	P��~�;�}�U�6���V��}%,��ƽ�E��>��k	��H�I�cTգ���MJ:�����]��:�{�D�21��+�>��F��7��@__�k���o��Cv3G�6^J��b����(�m�	��\�}��`=��$�%�`k�޽�\�V�O����t����g8�&��*�����|Nݎ��R!��@P�֩�C�(%��8Im����{�������9s����懲�� K*�����N:{�,C�er���ݙ�9��#�Z��vb����f��e)K�x�f͞m�i�K#-�s�OҾ�E�Mٲ�X5<����
y0ps�
!<�4��%��'�ۢ�+1�+R4���M��Vૅ*{+2�H)�^Zy�� i��O�n�5�1��7U�c�$��'���q�}��o&Ŏ��(E�4���r2=FE���I'�����f����1����m�7�����ʱ/<a���ʄ�l��� 7�a��ݻ+1��H���?4�/��nt.���$%�W �:
��&ܓzB�*�ƍINU���'�j�@oM�o�r�����`�@e�ص�JI`�Q���f�Z-�tH�b���E
A��f�R�n]Զ�������'����Ӭ'ћyuW�7�����=����+�<�O�:��{Zr?�T��z� �b"&Z�D5�MZH*��(*@W�Z�.UJ�K��Ⱥ����*��+}�\���j�OH�#�?�M7j����-�@e�+���Kd����^n���=ٶ>��x��b�����܏�ce�l8�Qfm��p:S#���?B,�بh�>k���cZ�%ڪ��/��Q-��˭�Qo*�M�i��x��d��)k**O$��L L���9��D���m�i��y��=�xT��Y7O�i]k��Ӻ�U-�Y��#�%k#w�R4hF��u,SHR�<4T骡��`ii�d���?���q�.������-�b��]R��$r,���&<��`o?����Si�bA.��0�.Z�7�ݛ|S� ��y׬���w!��u��?��H�l؊��4R����V�j,[���<���z���>/bM�����"�����]�F��\����z��53���,��<�(,k�sN�)/
}{uY�#�t�8���}�^�#;K��ϢF2Ʊ2��=�Y٥��Icy��G�?߬�G���D{�H8�Rk�I��B!(q��@K|������
��F�a�Z���k��t�	2��!bǂ�!!!�Fj���~L�[`��\�[*��L��޽�e{�f?�1��`�"t̓ �o�
cΜ1�֗$��5�'��jvE#����!C,B֠Z��t��JO��[���6�k��Cz{��ȭp��3� ]�I�Ԩ���U������u�IJ,e�;�6UJ�<�����������麊}��4=�ٳ�y�v}�������^iX����zra�%.��%�KVQL��Mz��&lJJ��v;������=�m��T�{v��d�b�Qf��'�t� <�I䡋ߡ$x���f߾��r��a6���X��1���e���!w��#x�~�gϮyLVw�e��\L���ADģ������m3I����ϛB�,����x�b�#?�E4 ��L8IFL�~w��!�@h���O�C� �T{ǒ��T�Vtc[0 M�Vۏ'�%^�B��߄���/�����r`v3�3�:$�ԃ?ju�d��q��f)�a�\��e70
7�k���5g,��.�k����b�"�~0�!��J4QiM$�f�BY�c��zOL>2�(^"�-KrR�&��
�~]��x���ݮ��f�WCF�5՜Ąغ/���-�K��dW���~3Q���V:��xEr�&�92 j�a�GI<��l�Ʈ%�w��;�P�u�7O���D.&��X�^�@*55��@�t�.�l2�l�0ϯw.��;�SLb�.��f�9plF��z�X�)��"4�:�"7��y�i��6-�֋X%+�v<����Ԇ��0$��оqK�t�Ǔ}�F&-"L�r-`�tGI��r�"2�2s����Hev�k�-N`1��??B_IX(U�6�#�ut�+�m�N��Çk
"�n�&c��d�.V��b�/���OΤ���HXWO�6�9ґ�L�4���)�՝���G
Tȅ���(&;�cX6����mi���_6���%��z��Súo�Dx05?�!v�Q�^^#�K	l�ϖ!E�J~����|�����>��+l�^(%ِs3-M�$s�����c��Q��e�2;XS0�hW"���9o ��-�g����v$j���E� ��L=��I�$ytV�Eg�{g��{�����c���\���TT,���ՌR|CA�����PVV�5�V���v���K?�P�Q����#���$]z�F�RNlH��z����ׯنhW�w�g���v~�
g��K��Z :��P6�ȵn-�q�/�V	��2��7ƏQA�7��C5=�Z�ZQ�i7��ΝX$�kR����A���g�)�lVV�Fk�`Q����������Rp��;���,_�+�2?lΩ����1���I�K���VI�n�ryLe'��RS����nN�����1����)\g1E�q֥�5�1'����f�����d����z�N�.�z�(&W^���YmA3���`A��0oq�'���g�7~�

�!�t������`�/���B�!`�v����h���$w,b�jZ� ����[��ʽ��`�9X.W�:��������k}�ÖR~� ���ٳr	 ����*(۶a�ݽe�3��xP��YܷT[��<�K�7�b�囅����E�4�w²gUq����.8��Hw%Eq��9K��ˈ�C��@b�0�I�0g*M��0��D�A ���I8	*!�W�! *��<��)?�#A�19r�`gŅE���&Fr�loL��@R��"bVE�X �w���.l�����WL��,�e@��Ç�5���;�O�s{�4����&9d�*��#
�*�Gfѐnt0�;�^��J�,�NM�,RS(�}�L���_1Iz1�?Xh�s(O��}O[E0װ�����(]I����E�3Q�@�$���z
iW�XaA���
��p��\聶I���� (V���k��������ne&1/�h#�E�%Pfm��>),B�B�7� C,�3�<J�I��vp���C�5P���W�Ա���I�&x&ҋN��]��&��-m�
��L)0���m���x�a+Wz͒��9I��SPTl�����z���e����mq�=Sp�x�nl�"=�,�^r�yֽ u�	֠@؆?ƓےGf�:�� ��N�'�����Vҫ�m��E�&����~D$Ņ,�`h8�k��鎍z�s9� c����o/]�,��Q��a�dq��<�_|ӦM�
����?Ùs����KD�cg��i>��+�G��8�ē����d~���|��1G���z��A~�U+�n�v�=Xk�D��O�5d�J�jZL�/����g���H�<x�!��V�Ay:R>D��#�ę���
��� �����)GV�|��1k��x+0�3�Y�E�d�r� nҠ�M�3�P�v�,�6�~�J1x��d�Q��]����v�!*`�⍛���v�H��A�BW��A��3,���9����b�
Zڻ[
0SEt��cԓ���I�Gq��;ßQp.**�<������[�%���7��ߍ�Da��Vf����.j�� ��O-�қ��d a��35E���:Mr�5m A�EޭO����
�Q���u����,h�2+���I2����f ��lr��0_I1�­[���G�:�#�������Bp�3II�~}>��`�#��$����J�B��N�?Հ0�q\^n�Y\Nwwڍ�H�G�uנ�������	�<�Kwu�p��ȉ�/�xρ a�=�T�	BEH���j` �d��u4��~'0���˲岏n�KI�6���E��������1rp�M�jÒ6G����k�/��ت��O�ľ;�%F����w�$���1z*v�a9�H����ML�j��?D��	�IA6�{S�w�"�@��Q�.���s^�֤�������E.pє��mg�^@���f �ȱ��(��� ���8��q%|
�������O||t����K��8�DZ<u�V�A �5D��sv�� m����]�鶜���+BjfI��CVhxh��H���%K�T�gvY���$W�I��8�i>h�Zr?i�@�v���>q.�i�4����?mC0N8|�\u�:z�d!��nٳG�j��( �`�s����U��c�b`P�`k�Zg̹���Ř����`���Pd�Z|}��ʐu�˝3f�>���~'��d��l�}6�Hv�an���J�MR�g�ӧqٷcx��ܼ9y����"�����g��L$���d��(�1�q�+�&�n]2�p��� Bv�l�@���yW�3������Z/��(���������j|��c���0��{G��l�7l�Ԓ�AЏ�����0<Qş�/]����臺�H��������,�.���.�;����㬈l���L+p6Z��6,6�Ԝ=��YZ��AD��L���I��xAW���:��7w�mS,���E�������C�5T���{�"�{#3����׹���.B������>���)�i�2��wFj�� H��=��pN��̢�2gP��jY!A�ޡ�$3Ӝ�ک��p$����@�͛~��=�y������R��J�H���Ѭ��5�U������GU�e��p�x�k`�{:]C�� u�q�k��X��?`�߿�9���zO>��`#WQ�z�܃lש��Q�ƛ�yјѥ^�%eЍ�_�Pq\ ]�q����e2<kaxT/~,NH%+�z�Ǭ����P>�Jx�H��-�m:#B�U/2�?I���|�R���&�D:�R�ot���ML��ne��O����E�Ŭ�3�2,��7d: k����1gP�S(���
�ᘡ�]q?b��!�2th.'�|~z&�P�GT�oз��ĠH�>���n�9l?�~���!��k�P����k0wŎa�I�F�h���=��V��İG4
e}>i=� �b��xH(d-6��,���A	�J+fU�*/guh.:L&�i�� ^�籌��g�py�5��a1���D�W_!��T���/�S?�I�C�n���_z!���4_r!��ev�3�����U�95d��Jd �N?'m� ��������z��"��@5=��m�F&o����1�ã�m��G��W��o6Ud-Q4�/U�0l������!�~/,`'����@.�e.;����诋7���f 1a���z���R{��0��~��� ��@̚Y��_�Zf��T�F��&6���
�*�>O��)�����+b����l�#kw�H�b�i��7�� f�lqh��!L��dY���Ӹ|+^&|�>A�%CyK!���=�+�I�"����Yb���5',r�s���#�Y���	8:������0{֬Y&*ƚh���|�݇�qM��	p��8��!6$J~a���O��Tƛ��Z
��Q�Z`�z j�'�|0���/����:�����ǩe��w���YN� �h��u�5��]�;D��o���~ӿ+UBD��<�dI������"CQ�d�#�cI�_$�d`� )!���i^$������F�T����ȫW��j��H���7V=3s��4vmwY�1)$Vx0�i�B�x��� ���	�C��[^�@v�ih,�zzQ/)���~�[�@��"�v�Ky�J�Wc�{�ߵ��<�_g�����09[�z�ѵjV��Ua{�����V��߳�Á���2\�K��y��O��'7�-(H�'m�y�ʕ��	˨���Ow�
#j_S�1!�*�`ň���@�y ��˅��I�_�!ʝ��f�:::D�"B������2�&v��|8dB!�||���_�h\;Ly�^!�k�����ZH#|LF�Ζ�'��:/� RF��{6�y���l�#��Ӊ�$V�6-�2?�4�����ˠ�JQp�̧��SM�6���P�YXf�x;�t#��(J���ЄFjFv����r�
�CS:6H6��@�ƥ{,��QftѲ�<�s�T$��U�]%�%�v�K�_F��j���L2��|�t@��_���#|v#ˉ��/p����8�N��]8�D�)0���a��у��Z�-btn�r�&��0/��2hLYdˎM���8S�M�Y�]�H�V@V��(C�=���������?0Hr�n�[(?s��J}U~IϤx����㊯Y��OŦI���Y��}=>��e�O�lTCV�b�E[2�����~%o�V!e����=�{"�լVC�dT� RȾ��?15u��=��7������܃
���wz��G�M"�Ӧ��%��uho�9���"������߇�g;v��Z��V5�hѢ�ۗ4�
 ��v&��ǆ������2gk��2�H�t���X���ɋ�0X�m9:�xs�#����'N�Ṅr����3�r�;���s�����״�{o8k:��k7�M�$ت�����'�g����׋���'�>�*� ��e�%_l
:����	�pJ}.�-:1���J�.��V����?�\e ;�ᤢ��F��)q+ޓ�ֽ@�9��߻!�mݓ�e/�O:wz�K�8�]7�m��w�c�y�\�{�wc�7w��8���v��ó�=��@�7K��˯D���<#�+$�vHC1�l��J���x�ȳ���-�(8�,'�e��z}E�4;/٩ ���OJi�n���`���h�ᒑ/�y���%������Kٺa����/�stT�ⴆ��Y��G��!Fg��uO����Js+��My\VH;g�&�[K���I�<}+=,�5
�v�xc`�(����/�ۼ�IAA�uw�5r�'����EtՄ����l��UC�Z��笐� k��Q�w�c����O�W��8R��㻓Lr���>�R������ƘԶu=��bb��`�]�X�0�;Wu�x�/���;��5I	]�z�d3;�*���ù��ŵuu��-0�G�k�_��'�8{{+���n��ƽ��`�W��W_������_[I��C�h�u�a�Z%u�c����li�@f-�~BRfE�(:zA�<]��O�i�{?k�a��1�L̛�;o���{�7mI#,�D�x��0	�E�5N��u��ƞ��ᛏy�"/#z7�������f����*�z�����Ԕ,F����IRyi�X-�����G|�f�5+�������������6KXL��Il���WW�y��\\d7m�Dt�$b�	z%#����䇗��,	�a�h���?�~>��(-�����j�h�2S���%Ad��t���
 ��ռ<W1��Ax>1-��,M��x���Vs�R7��5��6�%[�M[�z��\t�H	��&��u_"`�}�YI-W�Bo�]��b��g�����S=�����^�p��4w7�ޕ#:��#��U[���E�o^�!a7�lo�]����kq�w�.� �P�i��b1��������S�G�,! b���]�TB���a�/1;�I5��?������X^*/M�T���_�: ����,��Dk��`��$''c|#d�GN8F�*K��N{��I�r��)#6!n�4�����rr[��d�O<�;&�������ʏ�?w��r����5�gtd�g��h���uc<�P5��у�)x��_O� ����D��"QdAx���E����"�EY%x)�� ���4!�;QCB�KҤe�PU�7�2f�k�..�ml"��q��GG�)�?�`#�d'�U�5�������b��a��1<ޣuSB�u� ��ȗ��l���fkG�k�!�΁1���y���)e{���|v�w��XN8���a����_�O������e�`yֹo⿀���=k�����3GǍx�?��<����{�%�RQ�J�,�d	�B���H	%�($�v����XZl%	C#�؎�)�M*�/!{������i�����μ����>�}-�ϵ����;�파�l�_tjz�3		�{;-^��P����.}|�4T�Y�oߞ�Xએc_�Z,T�b#0i�R>�4͊�2���k
ހ��:�j*���O�:���H60�WT�<Ob
6-��q��RŶ�c��T�!s����{�c����6.�3��hIc��y�lΞs�'��'�-�?1��&�$>,�b��NAI���Y�Ǟ�=��D��k`^T�Q�S�LV&������n���'<�+�m�O_����\Bx[֯G�q_b��p�ڍ�/����'��-��`�4�Qgz<ed�m���ȃBFFܪ��*j�M���*�EsN�yT%���-µ��=I�S�}O? c]���4iۏ��ˋ{��"N��*;�93�-:��⩘��L� ���'�����N&%r�:��~��SI�8m�k�2���8Q�3��p��5u^j8
 .�K���I����Y�kh������v�.y�l�R�y��Q��s�:B_��)hj��@ss�R)M�+��U�%��e���ˏ9D�M���>bX��z�"-�Æ?ǅ�(Ql5ut���0MMM@�q�(Y �����}�)<3@���N'���7��L��q:��yG%����U�n�w`S�5L�:�w~�����? �w�p���L���S���+�1��q�l�W��+������	 ��$�#��Q�yyR�P��[��E9�^�ش9�1�����_A7�[���ӂL2P}�
ǃ ��H��u
WAA�OMIq?�L-=>�lߢ5
�$xC@?��َ���`�V�?&����-���iEQ����mC¥���g�W=k�d�ԓ� O�&n\��rh%�&�O9�5#����.�zo��]I�eH&{Y)�&��B��7Q���>����*O�% C��o$x���\�cP�.�I��DFr�i���G�~_*]T\�{�^�3P�����E2%�;�Nd��c��Kfpل^[f��p���0^�21�/��7�k1�tb�x-p�4�
ĩ�=\y����^�U����QT�,�v=b��|�z��.�tF�ˬ��r>}���@���Cû/���ׯgIM ��0&��|����
X��ٽ��󌚦��O����3/�r�=�0b�;J��m� �S�mv��z �,�h�,����3u�}�@�a$����x�;f���t���Z_��
w컟�j1���|)��s� @J5Bw$��Ş6К�Fj�o���U��e�%���o��[aN���b/�C`��	`^+��d��ķBO�&�K�k�1(C��,K�K<^��+rT`0�&7u=%8d��~с�}����S'��`��$�_fq^�}c0,=��k"�Ï8;�<IYp�W���x��b�-�XY-CM_j!�}H��6p��4/X�Xxp�z�9��]��cV�m��d8ȫW��L�)�~}���bg{��������M[D���&
�/���o{���jc��t��������eO���|0  �1����3�ѓ��� Qp#��E�$:��{�z�9��F�:(*���~��*p�6C.�����
�֭�+�#��'�0ڇ��Ÿ�p������ݚ�`p��w��IQ�1��[Z��y�'+�P
�"�0�}kTT怯
טҧO.u8a�J����bD����<�:�:���}0j���󫸷ӗ��z� _G�l_�3Z�H�	H!���"Eo�7o��1��:�{kc}�����$?xI�^��-Z{�M���>�������� ���M/�b���,�D4�������^�"���z���$
-r���P�����B��_x�b�x��`��� 1:�m�����UM/�,z��G3�;�	�k���S���W&�uC����1�fR�!�G,-e�͛G���L�(�������� ?�r0?�Un���%\711��6�b��	��Z��Gņ�kj_?�h�j���JL")�a�G�)RR�I��^�b����\?����NI�,��Դ�\S"������ĕ����ElW,� �{�^@V.���Uf��m:� ��֏b�>�a��$�u��&?�
��o,��UZJ3��*c��j�ʿ�d����G��d�|�wW�C(	&�-Y�����j�`L�9�j8>&��w~*Q!48�e�pz�+.Cw p4�e� �hİ���U$|.{Զ&~� �q_����>kҠ����&�vyU���rZ	�fkk�VC��'`aZ�M��D���Vp���e�B"�rwVu�It��N�Eo�9�_���J�\��r��P�����E�UThŋ;��>�:����?���O.޸}{{w蕮.Ѡ�ݑa�[�𔻟�IQ2�����=o�@˛z�����Π��;����zX,���wZ�-����`�H<�{��p)�Ɵ�Wq~7E5��s�Aڎ�S��������J�x�KTu�:M�0��l�δ��8��!�r���I
�s�,5���װ-V���:H[���k`[�Em��ح+��1�ԏ�( \���}�n���/��Я�i��������v�ewW�:XSI�M33�4�s�&o%�k�{�R����A}0�d䰒���5:��d�1�D�-��~�S35up	1F��Z�'@V�L���S���ӧY^^��S^^�#�������8��Ą`�˥��[o-��uY�=��?�"M|Zh��Ww?��«�=�}��7sm�����vT���B��G���	o.�|+��w�\������:� ,`݀�n~�oD�W��H����@2�bej2�Lђꖖ��� �Ck��ᔮ�kԶ���']϶�<[�a[��7n\�~��]�O�����jM,J�L&ֻ92�u���4r�5St�|�7Ԡ���7�LQ�=��B���g��ה�XV9���A�Y^��x��iL�9���0�BǄt�2�Tv}�]y���x���V+L���9 r  �☪�"P�G�m1��ͬ����9w���E��y�&ӚJ�/�`^�Dh�jp�d[�B��I{ߨ�K��
�� �a���N��ЩW��d8�f�3+��'���]�����|���h�j��H�~ݏ��a�o{�S6w��CB��:�u <$v�˲������&P��a]Ou��/?>[�.�p��5��
`�O���P�Ԅ�1��sմ��w&\W玾f%�lڸ_.v:��M>��4��d��+��,���SRR�� �񂂂H�=��=\$P�I�B�;$�]'&h$��R��Dg��1+��@�'�6�i}�9�T	�-4>��~���T�����r��GˢqL#װ�Ӫ�w۰�<*��o(l@sϖ~T�I�f�FRg���^m.�c�:�_eBƃuV���4���⳹���ܭ�j�Eɬ��9���]A#�+�W<���[�ڮ{M�����i�n��C��?
7���(V�9Rl���S�{��W�)�u�b�b�����R��A������S����7��U7
��B>�����;%�庁�e���qJ@`���1 �������m��n�oL���6b�>4j}DAP�)��{3�>��2\�L�a�d,�kp|��@���"�`͎0J��8,�\���r&F;'�:�E���YGW�H���d�\���g���(�oh�i7�`��G���]>�y�^l���My�:m��}�R�]$?�E���&�N�f�!��/�0�{�T����u̍�j�9��W�/�9�i_(�}����k�8	��m�'�t�b6�]K�<��qY��`�ߣ��hDJE$��h����uj'շO}��~�u��ӧ�+;��W�y��N�v&�A��3��`W�-�q�P[.�_<çi
bK�|p�U��g�� ��
�xLS����a!ӭL�����j��>�t�8�F--��7gh���L@Os��_��(���"��$��PRR���	v�b���P�G�UUm8�khq�`..�Y99��g�-I��v޿��"Z�����iz�IY�e�8���Q���7,A}8� LF��Q!�]�M����t�%q9K��(?���ogj��z�qW�9=�|�M��J5aS�Ś7>�ҟAB���ve� `�%w>Nᨂ?-�����l�� �L��vS�h�b�o�R��FH�N���7�m�;�@�͠{��LJt��+dee�LT}Hܼ!M�׼0N�[8��ӾJ�4�ܟXH���,���/�����KHB�~�؅�q{�͊�ϟɔC��栦��>��K+�ե�Ki=���Ϭ����V���[U�-���(a���k)�P*��d��	��� �D���'cl@:�����<	a���x��١'თ��n�3|n"魤f4� ���V�]F�a���ڤ��Y�K ���̫������8w��yդ�3�l�����.�]5��R{�����u�G��� gB.I�I�M�,�f����:F�a\u�O��x۠燝����l�fe���ضxtc�gϊ&�+]g`q�}�P�� K�
tSS���ik�H�1��sKf�oQ}O��"�L��yyR�d�Y��򝸷k�2�xh4��mNe�-���w��� ��w��t��#�����M�����(��S����;��~����kky%��ō�j�����+Ǵ|�T�w{�r�\�5?����f̎�$B�����nV�'�o�(��o��{��|k���
bP8o���4�/(����r/xi�#�E���=U��}��9����}kk���M�xb������4�K��jo��pݾYp2zN�.t�O�8�־Z��Z�#d���%z������Fߥ�/m2�A���R�VM��D'����K�U��&q^J�O�e�kj��;N�̳]qu#�	�ς�#�Y�yJ��h-ln&#����v�����:Ӯ�x�=����B�D��0�M����f5y^'2 ����t�uw�tun�N��/�|�k�g~=E]	]��K�Xi*~U 0Ұ���I�r�G�֋����f"��Ŏ�	Ɏv���[���=nPG�LQ�c�E�:��t�ع�?¹��س����Ԣ)�~���ɩF��S�jk��x3��_(T�G��ϛ>��q���'�Hb�z[�����H>����Q�o]X!�w�M�Uk�4��������k$Ϣ�d�z*@��<�?����rWWױu�Q�e��>}"Ѧ���J{W�������kX��[E��J1���1�5���)ސݓ���`8C:K�_yhX��:�^���g�(��3������I~+F21Gдcϊ�)m��e~S͑!�g�xa�H�h[��8ec#� Sv��
M���)��H;p���D����f���c`��~=i��6��]g!� 9V�UYX�u��tG Htv����CRd�nVq�o�`ծZ}��wZNø,S�C�s�h�-X\�;�}�_0���		8��z��悻F5b}Z	7��{�x�'���Iץ�>h��^�a1��::�9Y
l(����ck�a�7�$ô��Fa��*y�����%�Sb)Jle��1x|���5�3�E�.;�Hh���B�{2���f�TəX���%�O1�<*ڰ�8�0I{s >|@��@򼟲SS�i�
�WE|;-lϪG�T}����!5�qo���n]�hX�,�}1�=��m��f�Zl�)%r�2=���3g���W�g�^c������.� ���!x�2��7�>4��Y<˝��Z^��56!����F'e鐛?B�m�M��m�/�O�F����#���DL�O{�'Cݔ��M��?4C`E���ˇ�2�S{_�p4-���$!���zGUS+N?S,��%C_��g�:.8����h8C��uε�I�������ܯS�8�`y�Q���m@���(�#c�Y'�ӆZ-,��};��L��o�؉^1�Q8�H7��Ȯ��(��`�0��Z�t7E���[i��k���Z��Ԑئ/��{X��6X�3OM�0��C;iή���9p��R+vԞH~A඘�(�_��ǲ5+�7j�`#�����Ǐ[�`O����7gZ`�<6&�|:�x�ҁ~%��Z���5+�?CY=��W�����ly�]F��p&ݛ�y��G��ݸ��6x�)}2��U�j`<_�0��JQ`�v����L���a�Y���ж� ��I|Z�s����X1�T<��ƕ'0�;_��J�,Y��Z{3��g�����h�a�Hʒ�����������.@Y���չ�����g.�v6�mHt�r����I�H�17��j!����'3�~a<��0Cf5���hþ���Rg����^&}�b��ۊl�X���Y\!|�A�g�z����k�u
ooJ�p�w&mi�jk%#�bm�e���g�Xh�3�IM�����9�Fϰu�<���q+���B:�]X���	ceY�tt���`O\b���,�NW(.P3�;�9һ�U�ͺ�.m���Q����Z@�:s!�;��1H�}M��Y,k/(v�ZE]/�g�l,��=	|���d+���C.ag+A3̒���8W��JC 4C�蹍�L���pޫW>od���ޓ�t�S;S�C���t���ҡ��:JYg
�5�X�����7�X���n�d����F�����L�u��0iE���Dz�.�4~�����k�:N�jߐ���KKK'���k�}{O�p�;z~�>;�F0 �,��r��M(a2	��	���7���t�����X�1H:�ը���.z��C��h�s�����z,�dhE�70	Z�mC�e2_}�&�kj��'�+�te���I���Ų���{6���CdbhSt��ˮ��.l�h���^T�b^u���Cp��n��b�t~Ƀ��$-�`:����q����_����^>������(�,H��2�����/mą���ص&L����^�����M��n8g�π&��J�� kk����	�e����b��mړ#��[F���kv���7H�`g��4K�p��r:��U���\��af�)�ѣ9��=n����ƞU�GQ�9-n��Y1��;@/�*���ߵ��{�JuU�ltԝn�'(Nѻ/���TRs)���Aw	���z�x��-����A1�m�>�)��ډ>B �ձ�`�GF%��{RM�+��~�7���x��hMYX sJ���	�~-��]�Rq*�g�&{F-�W��pe��\��%R���P��q��������`�|��W9?�^ ��s�g�'e!Se�%9���������r��`���vڠsnKم�9J���t�V�k
�\�����S�	6#�C��>�Ν;�dE��[��&�S��Z�ksڋU��R�R�-�z�	K��
rw�nA�c��{Xvy��Sy��Nv�A�y�5�Ak���r���@��W~a�(r؜�/ ���y,F8ɜ<������	��NQ��í��e���X�I��z�����gM��ݣ��A��u������:M.��p?�{��89N��&9��T� O�Ux������z�Lܾ�-?Eс�a��`0�?<��,�#�1�k��/T���U���l�ࣕ����,�c0E��-�y�'P͑��-b!���z���=�i���1Xͼ4M���͋jp	N����̷"q��Y��8,!�D�h]�{X��1��`��g�'c�T�(N�@	~*/vqՕ
��K���0����0oȆpϫ-J�L��˒��X}�'p,�pM%�}���@��c�
�xZ�t���������#2�b��]��? wa�W�[ܫK�賜�����a��c����:'!\e���Uhk���!� ��}<��3b�_����Z�hA�F��j�H�H� ^�pĽ1̥߆�h���k6�[�^���օθ����S�x9��M���⦯�5��ŧ� O��cF?܎�u��%_jk� �AZjH���.â��k+A�t�O���9|x1=�mQ����m�~�3x�2;�9v��θ��K'q�=�0t�4(}���5��K1/�e������U���Y� ��ᤔ�V�B��B�6
 � ň�b?��V�h^xz/?�[Cs�
Ӑ�}��n媟>r���y�vd$�Kʽ�ڣ�BrnI�s�H��67p��pb��EN\��ULѠ:?يB�)J.Q�Ի7�g$tw��>��C���<��VQ������Yю���&!e��@N����9���:�14r0{�t�ݼ!�&�� �k�m�ɠ[� 	ش;q)�D���jH>��jv���oI:�Nٟ�����L�-�#���h<Y$y�k�V6���V��0*2�.�������>}�2}:R�U�v	����pܛ��w`�l.�^x�y����1L�w�W�j�ڢp�"jY��X����^�����"V&��w��W0�Ep��㣃�2Nz�Hna��-��+W>����LJÑ?啰���9�`��\Nya�Y����x��Gc��kN.<X#]!�W���#�#-8�+2 Y�Tc߿�Z�9@y�=��:�-:a�4̊1&.��.�t�y�c1�?����{(���?+;�������n�����p�Su��~:�>�����Gkc�sU�b*D�T��%�'�6ziU��Ґ�If�s�sO����8��p��M���.�pyŅ���	z�}t5;�ӧ�͎t�ͮ�=�w�0.�i����[7n��]lvT�$i�k����zZ�A�����-�a�܉��x|͂�8�q��q���B�'t�6%�d�����7,�e�4�9����[�{Cl�/b�J�ڪ�m'^�s�8Zy"�Xf��������Oυ���<E=��女^��������e�S�����2�i��̱�GE�b[�C�vJt?]���^�S8P�������˵�;-R�X�˜6���>�(�����5��+p-/r��#���ر���F�vr�]�	�$LcY(桑r��|�"E��emD��S*�n�6h�z���8�O?͊&,)�12���p�;u=������6��PT)͖)i�E�� � �;7��L��! 6���1�Le��t�8����E�W̝���;q�
2�>;.H��]�_U�Λ?�S�G�ꬂY��of�����W#ɢ��0��	�����n�ִ"���8�����e	���������-q� I$��`����"�ԗ&Yk�	yKN���Th�y~�Ʈ̺���Јqq���;�ҍ;̼�q ��w�]n�*j�Yn�us����u�6{�M���x��$���/E���ހ�x���ַ��&�f8c�!m3?ޘ$8c��¶������TM�W��t�$2�������X(]
C/���)��E��޻_j����� xæ�A��Hh	W��UQQQ�(�I�?H�ԧ:'���v])��݄(Є봃�}e��Z�[%�X"iڵ�h(���_k�L��~��1����� 9�T$����3�R���1�u��w�	H�]�)��C[k+�ϲWw`5z�^����p�83��>\0K�-=2�!;up]����3Ω����n��R�tT�+_ݵh��#ԍ�FU�G��%�^~�)���ʻ���p1C����-۷�p��v����h�߰�絲ky����g�$�n���AK
w7�XI�w\K��|����;Ĕ^z��Vr)�x����I=Z�Y#=11���n9Y������?�;n�ar2��D �m�^CC����x�]�	���U�S�%�P����tL���5��]J��˭Y�+����ua����:��6J76�XO]t<{3#��l���4>�*�*�p�����r�[���fF�r�.?Ni��즌�6�i1)�`,��i8��KX%���;�B/��م�td�<�����U��FZο�ľq��t��]�ɟ�:�q`͂�����b�K�EC�ǜѷ#J:�p�:^�8*z��퓹��@�[B��O����Nm[�y������1����ppv�_7K��[J�{$�$�#�I��i�MKJCAM����ss%1ddI�~|�l���cM$��ڗ��c���`�OV�N��z S�A~���s��q��%�2��P4�L�r�����&��q��R��A�W'2�J�	��5�g�q��G�qYF����.9ږ��8^C���l���O��l�'���m���\���y���h�o��t�Ҿ�x���O��t
�;���r�$~u'˂p)LMM�51v�*��*3'��S0�N}���}��}��в�._eJ�8nk��Rj�X�ܨ���%y�L�� ��˿{x�#ž_c�C����z����V��G�q*�8R�zZJ#��[� d�������?�{N�]��S�Lo���(����{�?X=�@`Ɓ�[���ϟǱ�ܱ/k�}�q��իW�8`�bρ+��d��ݡ�ۺ8r@�uҖ�z>�Ŭ/��Ξ};�%�,h����h�|i�A8T'�3,׀o<� �4����hL'��JDc�}EE���ю��5�pd*R>����TiO��3��ާ�%؂)�67�O��x�9(��N����#Z30�< �իW,��ڵ�,-xXNR��v��8���q�zyu��W�L�~̷��^��-E������!�_��ަ�b����d���%!�d� s�����|��b���A��oߜq6�23_I]���-� ��2l'��a�*�G���D���cJpF;S��=�X��.**��b�\��b2_�����T�}>;9Z��j�&�^$�����z_�L�T��9���`ƕ��A6�E�^��*jᰕ����<�V��Jjj7Ajn��H�n�h����2Fݤ����5��7�[$�h�w��V��68�����:��:�����L�{p@�E?W�)���yE��L+�dF�mI5��Rzw�{Q����H��ٷ��3�D�6������T k�|;z�����@���-�NJJ򮣸[P7�z��7b�8�c����~K��~�@w�U��/���,��3[9���[}jjz.�#�s�Ni�b�.�P-�83��#p�%�/��ˉ�� `gY�[�C����K���/��z�QkO��P�h�/ȟ1��n2�~&7*�L�m�pxW��L?8�k�%m��#����J��[�~]���?����>�<~�������[�n�K2��5���g�@��w��8nƸ͡���$c�:��}��5zɒA�o;�^��1��^Q� #��t
>�vq j���l$�c�Z�T�L�1@�Z�5^��40��3��

�B�:����e��D1\��U^s���s-{�	K�wHr���{w��T�+0��]��Ë����������IeI�aA,l�a˂��B�A�2&��i��������td��~�`��3��Z�����5�� 8�� I���M�\�ǜ&l��z;<��?9�w2 L.�*�\/�8���V&��rpi(���o����em7�V;»:��Z����$�U���ǅ^�'����I�T�ee�ee�������Kgs���m�7�aQ̾n*_E�Ӫ]�8��߆�4"Ӯ���顯;:N�x)�����J'@�?^ce���"?iӌ���O���x{K�������=֕�}�8MM��4���%�J7m�h�0uW
���#�*O�ŵ�'�)��.=8J�aq򾕠>�s͌O󳘧3�hq�z>\�*�-����a3
y�&��%tc�����@[Xq�Nb����c��^��OH�*1ȯ㰐�œ>�umm�c[=������1��TdL�7\T��X���� Ln/Y��EN'�t*�
��58�o⮌f��}�)�8�'��	SD%X��(3�bo?KZ�D�u�hȰm�6H�� �*;'�0L���3�[>��\��r����q*���֔:�\�~�O�Q>�a�{�ۨ�~�Prt�b�|��۪`�8�`�q ����l��F�y:
��{V��u�B�3�Q���?���hQ�ɼ:��CH�߾]=��`	+k:��)��G�~ၣ�DQ�矁�,sϾ���� ��7P����;v��*��+�5��0�GUE'�Ú�Vn���~?��xE&mN�H���NNxEFG�������u��b�'O~�d����y�����2z��U�����7��C�/��W��|G�¢�߹sQ�(���QޭkOl���(Au�EY��U���)X�,�-�Tf����+����Z+�(�밾�|'�%�4��v��o�ja�?��q&OK(֟f�������ᢐO.u[2 yƽ���g�&/�+��BT�}�9��ק8~{f :^6��Ъ���'<�u�X��9��#�R�3!�F��i���F'o�C����o�Ȅ�cӷ%e���Pfj� j���88(������c݋����p�X9b �my䌬0##���ϻ�;#�on^��zOOM�a���#x�Ŕ ��m��7�vw�Ŀ:�@=
t��I���
'�X�A�KHI��Y�G<�pG�Ͽω��.�����~ �^ެf�u������]���-A�|���-F�?}4��>��nDs���Z�_P��E��X����l㮶�
�}����W��@,4Pf�x���CT~-̿:j��;N�޶3ңX��0>WÝj�����R�����d�ߕPc�����_ [��FWrE'���KG�­H����Y� �bG H�H#�Z~���f'�� �K���_#xk`׽N"׌z�[e�Wv�eOf������̬�uܚ��| %j������{�cn�@��y�<�;��u��gz�Z��|��[9��)�`iu&w��S�R�W��u�ea����?k��K(�����h����������@m�Ži�̵tN��2�Z"���%O^��ђ������S��{��c��.f��<�M�(�W���r����>�4�D�(���[$��'�EM�d��g8�:Vb�g	��C�>���B8��xb�ϐ���-��c^ԈI�F�)J���Dft���rq�}
�)ډ'����7� �ĺ4��� C��u���
��8WLQ���Jۨ#Q®�.:!+_�($K�;�>������òX�|�7U��]'���K���w������Jw�Q�#̽/��KJ]��[�E��=4Z�}��\�K����gj4����t�3��il'wVIu�F�E5�)S6���	f���80���hx����G| �4M�r���C��njѻ�*������3Nh��u		����~i^��1 	���������ꅢ��GM�}�E�w��
}�{N��f,}w"�#����Y2Lـ/�?�;���J9V�M�`���7������1⹞#F�3��OLx#z'�[p�L��xv9k����� �2���#{�;�������ۓ�UN������k���Ԅ�^���Y��z�5x����.,�GC�0�e8m��tS��Z�j���8�.��W�_�m�w.'i\s�Ew�A����P�� gu�}��� )pDa0~����|�?�?����΄9�)�����JpF'2ge�1N#:�a��[#LC�S����C�[�n�<����F�~/;Gڰu7<b)|m��3w�1�-���G���$6'ȷ�b�(y�Z�1��nIU��l��: U��yYL�b�:x{G��q��o)�d��	�#y��HJR҉��;��@��?�G*.�/��X�v�\gIy��;�{n�/�}�v��Tg��l�Е�6�Km��B�Hߓg����!����f��|M�*�������6V��=��i;�O��V&3��19>X�G�	��Z�6�.�̚@%����5���0��iQʅp��-�6�ס����uO`�g��v:z;���%9,
2��%̓U�Ħ���쳗�������O_�?��qߺ|)h���^{���$ ��\7� ���X��-�ᎤT�� Njj`"�����Ӫ'<zt)��l�Ʊ�G4��@����]�6��?��$)��b^T¬F�'`8(�`�R�EC G���p�X�˫V�*^���Cz�#fO����	��~�$��M�~�x�~G8�m�:e�s0�EЎ\�{�& A��ch��:���/��:��7[��ؼ�i�GJHH<}��µ�l^�Ln�Çx^9g��Iƪ�N�Š����l��8�����FA�Lu­�p�#8/��������~�J�Es�'�Fo�-Xpf��f7
-�N�u��+�38���4�T�c�^hS��r3$$4�?QӶ2��9�A����*r�w~m��|�ڜ� �P�~cL ���@�p��7q�+����8Ʋ����z�����\�ѷ��� �XJ
v}z쟠Aeee��~�`���``z�u�S����1�RUJ��b��0��|�8�@��@�A�28�n-���6�U�����<id�7k��ԪC��m���ЕPU�qO)+>>G �!�s��hد�ٲILt\�������j���POYr���ф��P�%��0=}6�h�F����R����������or��=a�X�kƁ2�����Y��bǦb�h�[[I�/X�Q�)d������guD|��9n�f5&\φs��lߴ���;�}���,�^��p�NU5�����ck ���x�deK�q�:��]4ؕ��))5O�~c����){�����F��ƪ�p�����Mm���Im���g�gݿ�}�.�g��b�-I�6��A)�B��"n���9���U�J���~�Ժ�Gi��X]k�������I���m�[�k��π����вa�,@��p��֭�K0� a0���a4��K$n�^3��9�0�[e�E��Gt߰ ȷm'Sm�%��c��`��fQV}�t�����/Zyy�(�����`3�qZ������{�*u����������E�8�px	�f����]#��%6S-q�<��H\��qM�{�_���˗��������e֏�Wr���x��mt���o�V���<y�U��k��ݫ��Wi
��d�1>�ׁ�<N�4уq��J2��j�j�q�s�m��p��3 ���
�j��]ư�Yu����#2�נ�X����'�M�����+�����+h��9Go�!Ӫ�%>���«�|����׋ ES�lz�0_�,�)��ւ:��<��i��I�/cU"��3O��P!�LUgQgU*\;�D�����8(�}�c��` �a�`bt m�^��Zb ������׆B~x���3���' ��p�I8�b�o��n�R�g��z\3bյ�d�� �&��ٝ�!��7���:�j6�je�n
4����A�"i�O�>ӸW�{o���Q���N)��cbF0*k�5�e�ar��Y\ƙ�Q�3��i1}ހ3����
�����)A�2m�{W�,T=���~ȅs[e��-	�
g�r������4z�L�E��u04��a��߷�H��-��{6�pݘ+�3�_F����--V��<ê			�ŞQ�K�X=�}�a`��ϑ1�ʱ�6�+*��a�J��32p��5kB׋褁���������B�_�m$7�ӊ��C.��Ө���h�:��8�ʸB��t!>��Pnll,-#c�a��1i�
,�,��.����V��Y�3)��vqw_0�9}ZM&�m(���jė�XՂ�M���EeGw?�)_,5�r,��;���YY����`Xpɛ7o~J���E�!�ڀE{�Nװ�4.M�����yt����&���ׯ�H|3�J�B'f(�?�+�/_ƾiP%�N8�'&�Q>����j�h�!���߅����z)��2պ{����͔��bw��ުP�����`x�P�����q'��͛$7�}m�ӛ�+�I�%X?��2�b��_�_��8LLR�����tyo �p`ú��t��y6�<,}~]�o�~ʞ'�Y�W�&���9n��hѾ���Z�Ʊ��~X�vl��ȌzI))]����xy]�����J��Hc��`wعE'�T� �_�\�sZ踄=���yn�q������|���}��S��.���
{��bt�ኃ�x|�>�h���GM�ĥK��X4τs����H�E������b�m6�Ay^����S�d�j�Ǭ��?n��V@��@��6~��tq�;�~{�;�=��-%��`��C=(��NrXP��9�t �q��4#Y��͙�A��3�e���\=-���B�ދN;�Pv0y��/���H�YL;�^�a	��a�'x�P�ġ�G/T,�i[$t��$D:��6���~+��Q�A$C$u7���k?߶�sx�/�#P��E������8c�V�����d��3������wLS����'����#�_���A�0fd�ʜ��n� .wi�����q�ۀ���b$s���{L�q�ᑧ�1,�"+Y���2��_�P�6Ba�|�7��L��edd��6��(���T����MIV�+)�0���6���w�܉m�W	��y�y!��$0It��5,�


����'2:��z�<�+Bd����$�6��{����-�$��������ǆp(�����m�aa?>�j�s;m�O�+2�c_��Hg��H+q�bJׯ_7�=34xew觞�IlꚚ�{q��F)2��lvX�c�a�¶���`絈�O0K;��䍋I	��J(�_�`��^�__�tg�; ڀG�r�8��&�-�:��i �Vb���W�]�ۿNYY��8JB ���j q?��[1�k�0S�e��Ax�-r��k��1{�t�	�ncIEq�n���a�%:��|޼#t4���*O�h�}����E]�nu�w��/�H�2���=�I����s�M�X� ��_������;s�RY��$ QE�]��Laa=���%����<؋ӓ��������OT~7�qqq����&�����H���E.S�}�:o+�oL�`��z�g��!��G����鈱���B#��_c�;`)�o�A��d��l�n� ��2*90 �Q�2:�G^DKg�u���9K��d;�%��:�۰	dQh�|E3�L��LXK
W�<]�'OnO���$��-�����3@���x_��Ԫ��Q7�M�"�;*W�ph����*Dس`q��7�O�=J�5E���#'S5`�	B�K&.e�_�1KMh����̟X����N�2Q�;�b��T���/hŹ������h:
 ���r��������3V����bBpV0[0��ꓼ���ͤ��_o�������u1.ZM����4�'���<?x'��`�'Z*Ճ~{N���io��pb�~�����o]��:w�Y���U��M����r�IoȧlE\��w9:x2��ڇ�ꀶ���Oic��N�+!� �2���<c�Z�]���o涖F`jM�}�~��YQ2�õ��b/4�?|���{)^�Ng.Đ):��:
S�d�+����]�'�_}3m���!��K��@ܥ�������\���Ɲ��L�X�
X�Ftt0]��r(�����6�����v��GYD. �����X͊��S���f��5����'��G�wYYY\��9B�i6��p����S�e�6 �{עrr�����1��0�@�8yߡ%��택U$L[�=�%%U���1�x�A��}~��
B^K�;p�6H��N�v�����}Uݟ�#�2���g훪V:yr��� 9U�W2���Qw�O�e8�	�6>��'�%ʀ��ӗ
��M���� 
Hܙ���i�%�ռc��3/�0#s��� ����W �i@�߉R��`�Ձ��bR�P�l���¹@^0L�ܶ?{=N�$kxc�_����X&�Z�!!qݶһ-���1@���[��*�,����( io��w�X7K��*��H�Pg���V�f�^b�;w�t�;u��o ��"w�:y�ʼɉ1���^���2�bn�}b�o�֒ep.{u߬.���l+�� L45�(�5�Lix���W���P�v ��4<�	o I������<x��U�I��1�ǐ{�?ۥ�з~����
X��F��B��O�n� I"C�� 5�vu���,)-�����]8͏��ط�W�(��?C��x��[�c<?N]����j�cOm.h��3x9�@D�3���~�S���)9�^�I=
�X���_`ˣP�b-r�{�6�0�m��;�����Q�Z[���J�a���@-�6gQ�v�A0v��A's.n�2���/��;OO�@<��;g���wo����`ŝE+6M�S1wD����e��� ډ��_��_6��5�В�WE�e(4��zDOo�����e��]R�;#�J��
��c`r=����js�I����թ��C�hn��<x0 �h�F�Π�)a!*'����Dk���խ����/��v{e7'��{dٻw�pA�	-��2������v]X��kܫK$&�&GY�<���t��k2@8 ~�p��8|I�^eq��c|�)�klݔ�<��|� NK�^�N���72ZK�$����H6KՋ7�&ii�:�� ������9T�� .86##c{V��75=����eg�x���(�� �p����
���I�+ΐ��[x-g���k�jf��/��(F�60t�C�;`���1rF'�*΀�Hky^��q��ޜ�����~�`��O�}f���ܿ%Jž�;��6�"VqO�����0 ��]����W������7 5�I��3�}��ʗ����Im�{�b��D���:�-S�=g8!B�H �S�rln����� ���>hY!�`;eKWDlw���cc&�/�.�͑QQ8-�"8��m=�߰jWH�<˥Ǭc��~�����ʤfV���¹���j`�r_>��tyT���iKU2�y6[Kx22�W3R�e�{��=�^2����������kF�`��~��p��Zi�H���+�^}�F(Ԉ��?�p��t�]�y��[�$�G���w��$ϴ��S�[.�%X^��+���ݱ��t�D*(/1T@�p	;⨯�}}}�l`�G��}�����>|>l �m�;<r���t]���55g�����REG�<�K��/:�����e������&~2OB}cZ��b_�.�0�l�j��D[*P�H�j�4����k �D�r�t����5�.E���  f;F��_��R5t�2����%��SSKR�'����9#kqq�4M��(@m[��/5������!�(^ SGM���N.��cQn>��p �%D'3��a�ѣ9eǪw�f7$���k͵� b�����#k��)�XE��6��b7ɐ�Y� 1�!`W���"�M5f�x�������4Bx�M*�?t̕�G�>��M���)�;4��<���.�����F��Mg�Zk�Sb��ܙT{'��W�M�˯y��r_u�H�т6���v"��{- `�X A8�����&)e�D�8�8QBBBb%�-Y�7�[K��B�<�5kD+�T�VmP�`e��+�ފ�~5uP�k�y�+C��� |N��^tb"Oq%��o���#�3c��o{�v�b�M��#��J���G1�D�5@j���cU�<�ep\eM�/\�$�����9�"����~��qO3#��)���v�������y�T�YD�����\�ݸ��z�� �`�'�0�}6x�\(� ����"�] �p=1l.�������iW�	�8gT��SPWW�[e�=s��Z�ó@���ӽG���{�wQ�Xݎ^�R��M�:O�Վ���ؾ���;*ZZ��:�Y�f
=u�!�v���ЍanD�����~�X&��c�[PnC���q�m$뱙���O�bϼԼ��s]b��o�[y">��'h��|�}�y���m7փ
Q>������.a�Yܿ�h���㘄�)�[j����z�;x3Aݰ����w���i��q~�p�bl'��UD�X9��	zN��m��U�pec���Q�椭�s��T}��`�Uj*�aicS�&�����Lj:�5�ěr���+�ލ�_�ҕ��n���7S-O@��Ct~F̞��5��p�ue�h�g�ᙥh^��B�����G\|Q�:�{u�M�f)Ƒ�7�:����kI�����PM��O�/\��x`�kw7�~����>;4�FZ�p�d�����*�G�:��W��g��^���\��.��d穿=�>����h��dG���E&q���{�xRGކ�q)��%z ���JN��}��� ���3W���vLSZݯ��Q���Z\�-FQlG| �{r��ޡ�4�Io;i�7z�P��.g�-�Gl�Bj��*����n\Ê%����7o��?:�Ѽ� ��`�mU2�+��fԮaYܛzp
)�H��,�ɗF :�����4�I�G�c�|&�⍘����O{+bqo��.�Y�N������$m��~B����c?��q��]���A�8sN.�4؅\��$c<#-M�*,��f�� u}`I�J�l)��l��w��A1���&�~���N�ek�i��^0H���p�8I����h�s�����]�匚��X��ئ�����@(����$���RT(E)�XnDQ]EbJ�"K�,3RQ�V�f+�u%Ke�6�T��!"��e0�s�������~���3���y��>Vc6��s�ԩ�+V�*/f����j�C�h�L����j��'1츅��l^6��Y��ź�dP�C��^�GA����g���\T~Ն\�_��悗Fr��g�Zp�R����NxE.���`7
rL��}l8�#kw�����ҋA���s��]��e����(SC�M�~G��B���u(p��8WV%F�:�����c�®�p����d��q7��
��8��-]��}��d� ,�;��4�E��B2��(��}ͱ�Vu��j)��Z��M���@����N�O�_�/�bqͬ��k��6mڙ�Ctk�6�g;�@_uS���H���&7d�DJi�.�?o��]���a�H��廬�q~��ygE�>o�4��EL^�֕g8� P��h"���|"|iu��}�IM� ]8I�~�s��ɷf�X��-ܱ5�Z�>CF�Ri�xy^�7�R�KEV?���l�04���u��VDJ��Yl���u{g$1��h':�|AJ����s36�5,h1eׁ?�h����P3�YX�,X�L�CȾ��)(�SԢ��g��*�����e5ִc�b�B��I��52����I=i��}V�N���w�� (�öov�{#�+"6s���2˄ތPșE�s�l�ho��4��5�2���~����䕀���0�{�Y
��,v�G�J��<�Cf��`QUU*�y��y����U�t-u�|�a�Ѯ��JG� ��x�LW�׶[(��AZ��Һ�(
ҁ��C��|�f�i3��ff.!������O����"%4�)�o�5���@8ߦ�S���xº-p���%���y5]e��`y��:Xr54u�:v��eTX��'��+pBV.!G��6�[v���9��ȴ��}��}���ɀ]�=�*��~�\�d�������=�v��Ϟ�:�E�T�@��� ����`���/��S�{�&�#������u-��B�������Fܗk�~��)	�ƞ1��.A𽿲L��oq���o��[&Y�?�^����~4���'Q~�ʣ:s���������[Dfx*p�^??S�0imoo�GRk��X�$2�v������T�q��d��!ګ�l��a��8��u <�p�jϥ�����7�5�W�o[G������<�B6v��u�vsf��()2��u�����AQ:���O*|��p���w}��_�C��	XĊ�0�d!�w��
~!�]�<�����{cw?�����\�v��V6��;h7 E��X�m��w^�<Y>��^ǟ&�;&`���Xҁs��E�i���a����H�6e>CE˭���?���Ƭ�F�GXlػDN�am$qzBR�_��#��̒�����i�[�sɡ�n���]�׆�1Gx�q����Ǳ�l�5��2�S�=c��� m�C԰����`'*���kUZ���r�s�o�� �z�ӥB��0{�-���6���7��^���w� � �I�=$���x),��ɩ�-��~��!6�qrv~y�9%!p��ۈ��K�xϸ3b�d|��/�,��K	A=�㒘->0��q��qW��2#���	;��)p���+o�,�ߜ��6[O�ƀxq.a2�&.ɉ�:�LY�8��5�]7�s����X���l�Y;H��S_��D�Y�1�W�,jF���[����뚆��*��F���.�`�b������f�iii����;��d^������H�'?���a�ߧ��2�t`C�ۛr���f|�|�U�$�=�:r�Z��c�����؋cll���_J%3�~��'_��U g#���\J�ٺ�1Ž�o�X�j�ID�C��w+��[�$0�KO�C�k Y+8�z��%1���:#ѕs�������G�X�(v�M�{�U���m��O��(��c���NN8����?|�d�"5n�E-�\�H�w���b�W2�#[�݋������~p�ȃ�˻n�60v�l���i�d������9������}����^��U���H���$;�ʈĐ���D�L��;w�������g���9��M���h�n� -�m)�O�t����3ǖ66^��[K��o���}��.��A\��!��%6H�ԍ́�E^���~4!�`��Ffm���A~@�ۏݪ��~d�'�t>�\�-ZD/��p8�^�ϿYl�U��"��(��g���[����i���չ���n��:�p�9�Ղ�`P޽3������M���>74��8����������GQ�Dv<m�#yߵ�Mw��")�`�C�a�I��=��x6Ol�p SU{ǘ�˫ �@;0S�ׯ��Vp)/��_|ʣ�H+?�}�.,Y�%p�_/�D)��ь[��-�f��bɒ�N%Y�o�yd��ֵ"?5옏��S�M���h+F��X�ǹ����_NN� [1���݅R�ڀy4G���5���t�s�ی��0�Βo�t�Itzp 4�9{����A[�r��{��<�������~=@@�p��f�}����*G(p<74_�>|8�u�hq�Z�3�p3���M�� �ۆ����lC�@q]���Z�eh�-ԘKG�&�o��zc�5<�g�X����8;��(\>�[2�B!�>0��~o߾�Tў���.[�4A'N�O�2�>�Rc��ǟ#���m_V$��J���l}���?�$�8n�y������s/��d-5S��E��`'����������� �y�+:ޟe���M�p6UZ�n�������Lq��[���|����ly� �c L�J	�?�_F@��ѓG���`E	'�|�qC�]�N�5F�	�2,p���)���"�@=?�JhzȓǇCG�n��l�	�Q^橘���ƹ࿀�c�7�W^YY�k���`N����W�wX�p��H���tɞK%U�S��~�����-�2h�=���qrC������������7(�����%�0�|��Ƭ�י���V���<��Ht��G�n�N̑Qwk7@��\�۟���ԥ$�h��z�h��Ne*��5Jy�'3��n1=}��!"�D�oӎk�R>��>���N� �֢�4+�N�B.�)v#�%O�t���;5�5��ߎ��'�`��y����v�>�!K���USK������|���I�t��J{�����4A�qa��+���A�?��������w� �`�!?u����ZCG�8�MCҁ�3d��\�a��Wm�������UD������N�կ$t#&eJe���x�Й��"q�!���H�2X�g��QX�k߮"[%�����
.�Z�G�Y������I�o��!�]5��Z���7s}�$/��3vk5^g�7�Avl�OS@>̿��3O?��p q�݉�d���ί "�1s�7���P��=D*��p��Y3蠡� �@�(����~p㐶�|�ϙ��+����?vw��/y�=���zP&჻�"������������xn7IaԾ�:�|l�K��YΏ32��-��T��f�QE~a���C�$�%y&��	i�w��`#tП��٦�"����e3j���`���~8�o4�,�Am�q�g��gA>!� L��_,%��èWw��t���x��=��E����W���l��X��ۂ_�H���a�A����쬌�,V�O��p�eY�`�Ԇ�6��j.�`�Fq��~b�	�K�S�]�ۃ�F����t\��r��/Dk*�2�.
^S��ą��lt3`�1��FT�7FQ�����GE �~�����F[����sZ��_�6���R��K��|� 	����L�����I��t�����Bc5�o�nnn��L�ZLN]�����`�J�?�����p�r���j��d�]�c��4K��� �,)d�8禵��iADD�XN��8#*�Wg}�[��M�����ϟ?�%���|�5?i�� D8v�T?�c�/q�Ej4���Q��������XL�.�H=P�EB�4�ķ�ۻPjhs#༝8q�"�ߺ�f�'VF�s�0����	�}�C��2V.�s��&�s�w�>AQL�x|���1v��/����m�U�ƀ�� �p�o�	lr_C�����	�e������_9��`ظ�:�:!)�8�f����l@&�T����t���G���E���wUD���=�~�I��z��p$���M��v��mۓ%`\���0A��|��ݠ��Ц���ӊ����2m�'0m�^|��6�'''OV���`DcPO	l_Ӵ'B!�� �Ğ[o��dz˯�q�]�/y���C�׾�Hmn�� �i�<�8P_j��',u!�|2�x>0O=����iJR�5RZW
l,Y��R�.c�:M�8��4� ���-����\����8�����0k��!]¿�	u�ո�X���df7S�>G�ׯo��$���t�S��������[�	X���iM� ���e��T�9�UV�N_q��p{3ynn�w��`�be;���\��ەd�M|�
�f��퀵�y%�lN�|)�.�k z`i6�OGl�?a���Y��4�-�ROs���}�d��	��S�G���_p�;ܑY�WS>t{ܚ�_��)	ε\���N�ȘkfJF��`ִle6�V���[pԛ�v�������h%�0I����.�����c�$'č�o��#���R���s&���1Y�R�D-��WC6����ws��q��F�;���9��k�N��*�=W��[��`���w:����e�V�뗳Vd���cz�����[;��
Re�Ij� �EWϳ	�}��⡄@|y�k`�	���t�K�ᯢ�y���(���	�ȫ����� ;���܋�= l�R���l�\�R tu��{����J\����B�_�O����O�W��{�M�,�Y�Y�(�^)�>u�(�b�`�)��{��H���԰B�$,�
����_����ɛ���Gq�	�ӧ$t�''澡���r��lQQ�Ħ�؂�u{�@5����H}�c)f	�d�ݥ�97�ی�%]��wk�����G\�9��D�����;��
[qM� <U �-`��˫`���(����]�%�U55A<��x�ĸ��k៱/'�\�$�+���@��8v����qW`����63]F��e<��Z"q�Ъ����\�o&�q�g���v��#��)
Y�-r�`��}.���V����H��`%��lq���!�͸�,�驣:�:3�X���s�!r.�����4��q���t��M�� d���T���-�T�a������z� ����ACCn�o�n�O�D��͛��ۗ����Ζ�(+����sj�gO4��e���!˴�ط����@��e�c�'�<�a�����7�y��=}���6�k1���am�֭��U���9�}�C��P"�ؗ.�͒'u��[�<7�Kn����_��}d�1��߹����:��	�́ ����M��-�_�B"�2�����@mr�[}�q�-v�h�gF���@t � ��'���&�w��MӅ_�e��<�k0��\^ᷞ��[���排q�(��-�vt�_�ǲA�[@���B�5����;1���%����i�8���(霫��h3�i��� �v�t�z2D��L��7vO��u�������v��h���ocr�@��ͪď�O�
q~cr�-�����Zn}F��y����X���0r�z��X���By�;ǚ����cI��w+v����l~�h5�����%F�Kc��7	�>La�	��}MHj��~323Q�?�.�f�Vu�LL���f��hc^�����V�Zަ��]~���ԭ�O���� �[���3	�ov=Ԁ͓�8�[�js�]�e��s8R�����1�#�82p}Sf[<���}�9�u���B�ǣ mx��q���*
��<�2Np3'�S���݉6�� 0�]�Ey�/s�K;�lS\�(�|��:�t\�˦�n��.Y�k:z�FT�����~[���[&A�)�lO��s��S�8wȭ����%t)�6N9o��>)r����|�'����!C�/ߎP^QZ�r�cu��G�u�K������J�xYd���oAO,����v��u�;�1��߈����ns3S���t�4?����c�a��j��O��{�f�����I,�#��� ���̽���=<z����G���f����m�����mlN:ͨw}�%�;��1
�~�>h{E˻�g1��ה]�{�UD���cg*�yq�?��E��E�y)�-��mj�n����<�!�>g�gvlI`W�?���%v�Q`�m��2m�Qx�MM�����Z��l�@�d?��Ƽ�w��Kd�̝G��f`X�np�|��a�_�rF���]P5̢�G%;c������红�Nn����Yc�nP͕��᫷+ѿ�)F�H�m0�O�6�ʊ|�����'�|v�t�%�$4���X�U�y) �^���\&gZ�i�'�p���>&	�(Ԍ`����CP�S�V�Ɋ���1,�]87j��4���283�	��/�C&��e�(��0k�Rl]�U�i�i8IN���5_�=��"�۷ǲyjCUp(��N�w�V�34#�����KLJ|������"�3��{l\��(<��H��8o�o�~;+�jPƾ�i$�a�O���>���r�r�PG9oP���^.f>˚ ��I?�i��t��t�;HW�1�D�@6�Ug6S�Ź�IQ��n�:�}L���/-��D�����Nn�!{%y��Ht���'�U7��_����y��͎e�yF9�g~x���aꏍ��\�f ��ZXj�>@�z;�6y�����#���[,E+�k����qיS��qGc|������%���a�xM��L��bu�6=�k�0q���2yD�?��p�x�&���r��i.�"��fGYE�n��l��pEK%S��!H;��������e]j��2�E������)��ڒ�P��l7�x�UCThɮ8�\`V��WT�w�e��m3n���t���������W�m�q�[(���qM�m&����y���E �a���]׬p�ytS�0�������@8"���:Vch�� 5��މ��+e���S���.)X!�v�%QPFn�\f�!I�`{��緑�bP�$=�J9G��ŧ�������Ꮹ�CnF�����%���
��N����}h��E =%R���p�3,�&W��>/�#�5�N�pX��N��8�lq�"K,ս��f9Ь����K�$�y��d~��/�zC�]����T'躜7ϊ�@n�rc?��� |+,�dru֫���a�����n0�W��ws���	�N��)�tA*&K�<9ܥ��tT�����F�h�0���� �mm0��|�X� ��{~ب<&me�F�?��%E=���ʹL��{�u>Aw���<�[X*b*u�C��x�7�]�ɾ�;~yh:o� �$�ã0?D ��s��fu�OG|]����8b��1sW�a+��D��0��/	�7�:�u�!��pm��ۮs=W�7�[�P��V��͎a�o���hnϸ��U4�L��{Qlȥ���W�飿��ոc��0�v�Q�}+�YQ�D���r����.]��j#��,J�ӛ��&w���b^�Ď�԰[AfB�j���������5t����%�`����Z�a����yD������Ħwٽ5���O�sN��6�#u4<��a�y��6y��%�+��	ųT�47���+�)¹^Ն�w�Ƿߵ�,($4�f�F|�H��L�3�:R��1Vow%��v�J�Y�@��
d���~h�n�ɕ��\g���4 l��#H�����8tk7NT�`jT��=�M�ҕT��u���dc|�^����dR<\��	�����*���:K�7�p����S&�� ����"�Q�0�a)��ig�iE�����J�`A���3�%�	����9oQ������Q�+��
m��k{>�.@=���z[�s�l�C�ds2q�y��H�A�nXhH�>%C��r@(�Ps{�s'�ۍ��M�`S��n�G�}$TE�["<
��-���͂=��#/<N������Dz�� )��k*��΂~FJj�YC���詴���#ɤLEg8�#dtf�Hs��O�3��L)��E�Ӻ���N2��ϩ��{
�sz���{�*�9F���Q��W	3o�E���$jd9��D=�>y��v#+���_^�@R�}K@d0�W9�;E喖��Q�68��D8��?ioi��w�à�G��I�
��p��h]ϘOG���� ~�Cpj�y�D>ԫ@�(��3U�0?AM���tJv|�x�h`v����g���&�����g�S�:��pP��@=�A��b~�@��k����]x+&�p ��$�yEΆʭQ�n&�� �[�7*^��*I�@�@5���$G�T�k�0�/ ӿ�������[6�	�ytdG3��Rݝ��.��.U�dbR�6=�M����#�aJ���+��L�[w�W�����\Dâb����q#f��W)5�l-@�14}���E��,��=���AOzE�.�!@�jy�6���X68ri��Ndf��_�k� p�(�k��������T�h�W���8oWH8\��U�\���ιѓ|��Lb6{ʶ'�����	��xm?s#�ma&�p��p���Y���3S#8�Ȉk�q�����Fѻd�� ��-#���zH1[q�&��Ν����R>]q�zo�94��Cl�)� L\���֏[Ey��H��3���Ē���I����p�B���9�_�{G�?�O�^����Ď����r���>Z@0����<�?S#sL�3��&3?������v�e���jKP���̎�����y�k9�^F��Z�=�+~�OYJL>�`��%����-0��)+�s����Y���O� ���t5{����� ���{/(VιxX0'E��ԓ����^����=~�Y�@,j��8mzq�ҭ�1��S$t�ćĶ��l0���lU�*�@^��C��?����0���+��(��A�Y�~1V�Qg�l4 �I����'�5��~������'N<80<��N�gN�RhM ��gC�=����P�4��E���0�G�2�q��g�ZٻfR�����55���z�{�GF�l�W���1&�Ns��Ůx�w�%9b[?v�5h�ں����e*�;5D��Q]�WR�����|�l��<���+�gA����Έ_R���8F7���7�4{X8�֐���q
��P�***�7� 
?�ݺ�M�ؗ��#�@_V�_f؃g
����[yX�B]�'�)}���ٝ���&.T��>(�X��F� ��ra��\?.�ゲ�狤~�LC�}@ݳo߾�֔��ס@�N��D2����caaaCÕJdgL=i���8wU����B�d�ܯk@~�6�x�/-��S�$��E�*�g�ޝ�oms��L��nΫ�&����%�E����y#q��C]!o�tKV�L{�/	;Η�P���"֠�5#����]oc��r�[.~��ϟ'~Ϳ���*�}��\�r���4���	ŀd�g��%���(>w�L��H*�%2щ_��ji��(�&���WR�!���|�{R�7�>/���Ј�Rp�˵	�fX�,��s��7#OA>�t˰��@-��9%5d��*9��}?��،�v����[d;}~�6�B;�Qf�Πv/���[Vnf�9;�Y0�� Uj�|P��<�ބs�8T���I���{����"��g���o�Ct�4�� �<w�0%0t����� ���y���J�����>��
��d��؈4����(y;2Ӛ\-,��g]	/���VGJ����o�Ayy9�I�u�073Հ^�<���ܼ�	 7K��
�_ث=�ݏ����R�{��YF�*��(����⃱�)� ?���s���uSp�6���/-�J9z�7�-��Xi��C�n5����;���vSO��M�n�:����lE������v��ث���]sh\l�8�L��R�K_~kE)�m�"8����Қ�p@��F��jEi�<ȱ2Xh���?n����sGf<ߑϛӯ��=��4��c���`x�#����2��[*��G�=��e\S��n�Y�v�b�0�p��e���������d�+(g�AP��aN(g��g����k�]�-e���v�&)\�̰k��A	�������v�ʉ��[�8���`m��T8��hP��g��M�,�d���"�8�C���eS���muLG+b$�a�^#y
�w�n�7�o>��֌�o� a�Aw����}����HX䣶�Z��v�e���^]��{#+�ʆ)d##>'��o>��O@-���K]��,�`=�`��l����1�b�OV�N^s�Y��lQɄ��SA�	�S��H���A�s#*c��b����ҰV������ȁ."��8�LE��S�F` km��46�p�s҆i�	M�>�	._�x|���T*�<.a��x�+�m3���5#'�O��e�IHP�"F/H�n��]��\j��ո�R�RGnB����*j)��s\;�xRmD�9��Ô�� �����i���`6p��<�*���w��0��[�gy�N�w��XY[_���� �;�R�8��r����y�u-l�"��ӆ�"3d�i�L�@EG[���{�ǝPգŪ���͈���U���pX�;=��:��ip�g����Gw�����F�X�$�[�,���)g�cV8�w��Q 3��*���UzI��#�%2��Ӆ�� �����(ոo�<�	�j�n��V�j[+��C׿����k�V��awk+�i+�0����׉́����t9��m�����G��wg��$�����O�?��]G]����ꦭ�aYYE[�K���7��=S��u�� َ�c��]U������o�����A�����|��l��H�v��;�+�N�{�m��wы�l��Rw��d�w�2|`B�L�����R#͹��Ԫ�*_~�g��UZl){������� ��
"=�K���7�Wb�	ЂC��0874��B���#��.���΋��ܺj��+�M�Z�jp6,�m���*��BW�[��c�a�#�;�����Y�Xn?׶xn5'�yC"}_�L�?��g�{���B��D˴����i�i�"�C�u�f��/f.��C��X \��>F�z�*�?7�<L���ǯ������@�Zf��S��\�?�4U\���Q�;�+���V�3�&�G��s��r�m�`a�A��j�̢��mb����Ю܊,�L�E���̩�4S*=� lÂ���7����N�u��T+f����UzmX�6|�`ƻ`����KK��*���<��U�畮��iٲeC_����Q���VFL�ҝ�w����T����4z��wpį���7~'~h�]��K�J1U~��B�9<����ZY�G��~=��c�Wv�Q��e/�sT<3������3c�#����X�p�}�7�궷���
Un��yl�Ve�Id3v��ΙQdv�+7�8j����:���&3<�k�b�|��W��-/�y�ϝۊ�7@�V�)7�s���Q���M�]g6�� $4s�R�EQ��	���?}�he�b�8�:������؊��~���AVk�?ZA��tgǛ��Y/����꺸�#����O�����q<��ڗV�f�z�Ӆc4l\��R"	�,`l<�z��奅hCS}�1<�'��԰��;�{sL�y�kBg"�n�;<��X������������f��u�����Y����9�J�8N<�
�2��h�T �xH�����_�箮p�d�:��@�t�������� �g7P*M��A�+���#U�������6��+9��̯�d[D;H0Ex��J� ���(�����3�U[[r�p$r�7>j77;�I6�D�9�/��B |�57�m�+Q4�g�|-+!�JQt��]p�>���s�|�i�g<<���Y��5���s^�:V�v���N,/�s;)�����>k��<J�[Q�k�����\ �?W4�Y.9��Ǐ��dWp��ؔ��K VR��rJ�u<A�F#��]�D/���(ӝ	ag
�ϗ�d�87�Q令�lk�i��X��c�1l���o�#��|���*���Ι����hp� ������z*�p������ѣ���p�'�>'E����, Wl�YՖ��훮�젤Ft��+:����;uloIST �*��]�T�*��ιgLD�1���+=�i�F���ɜ܉�s�����(6�g\��	�BThue`$���3l4� R��
I�����Qu���x�����c�G��5sԯ �0ۓ9y����p�K��#����-o�j�^S�����^�8{h*�:+P>�Z3AJ5l�G`��a�3�M��&ɑ�_����|ev��ƚ���,�o�����9�2CCCA�� $=p��<IuWl���޲��18� ~9��XOڸ�����˽A�?�|y!,Q��1L��?��ūб�똋��j,2:�!ٔK(�z	�����MWn�@<S����@	xo��k����/�T���������s�?�E-R�F?�d�J[	�*dS?�E??P417:I�eʭ_�Ì�������P��c��رf�<OLh¼��Imm���~~�n/�TQ�7/�,0�Q��f��yyx|�(.?���^��R����i��E0��&D�s
�c�4�/����4>�s��
,���X�T�M�����[d����c��gq��9yQEEڇ�}�e+�%̍��a�;,��榃�̐4�\á
W���|�~z̀���@�ã�R��Q���:���ƕ�~8���N����f��[�ɟW\�?[h}�VtpSe6&*ǜ:�`|^;�	�R_��1'�VG��M҇I��1��;�d�'q�<9�K��>L+��PGE�E�p�����5>u�n^��o~�Ja�;_�U��T\�5�.��l7Sn�{�j�N�u�ж%c�[\�$d�ǉ���uD�}�QکE����b��7c�U��k}}���^ᣑ�7�d�&D���I%�S�훹�����ok�t
`]$_Y��ġgtd#܈�
�5~~l��Ʀ�x	ź�X?����j�����`�_�τ"����;����6�������Ȉ쎀)-���4�C�2O-%�����g_Xet�5 �lJ|�J���q���-�m9�n[�O\\D���4�r
��hA��-a����Q���?`�z�n���X35�Aw:�`��q���/�_p����y�Эx�c�z@�0�)�b�n�ֱ8S�GB"'��x��X%�Ɇ�b]����w�L���̅�������q�ހ%���l����/a"y��@�|X}�H�AB5*e�M�l�␥��N�e��t'�u���|.�^���DJ/]��Lۖls�o�ohh�E~��C6�ƝD�q����JN2 (�ã^�Ss�1hH���+i���L�5��������HJ���k���(F^�ə��2} ������	��a�w�$WS�F�U�t�x-O��O3��;&t�M��~�\6��D�����[�7����,�-�\���}�	���do\��22���N.�@��Aؑ|��:N��2+��*�Sx�&a��J|�P�M��� �)Z_466��#TZ9�a���㸗G�M�t�7��ʕ]>�	��w�T�Ut�x^kM��3����1���0?efjd���\��D��?��;}�j�����>�R1GF���N�یz��(�,�&��<B�
xC�U�* o�����d�kB�n���U{��������ޟ�ϖ�]1��b�D��H�4=r!����+x4�����=tl�&%%��]&���&��uY�ئ9m�IT����lj�O�<�J����{��KQ���tc������vPjcC����S��s��0Vؖ6�2͸����(�<�`^rr2>����ud���G_�"�t��}������"�.0����_�� ���>7z�E��b1��\��[�p×��;��%d��z�v}�+��	 rP��M����I^2�l���1�yNn�@�� ��d��No�x�:��2�gF~�i������g E�����hlX��� pUہ v�U>�cy��e`s�=�d�%�c~xx8ى�O�{�I�셁B�t<��G^`�40��o�0�p�+����ӕ��ыv��%�mu�!���r��d�X>�&�C� .^l�������i �	V66�;JC��C����c��c����@Atg(5-�Ɩ���:G�S�� ��D��l|<G6v�C,1�XűZ�t޴m<of��%�a rm(���<^�~���H�(V
?��τAҧ���]+�QUQ8�T^4,'Ɂ�@���m/Bw�.(XEb6�O&3nt&�脣=c��d]F��@�"�ʛݸw%�(����+�������9� �ް��T0�y�7b���>�)ҺT������N�n�yMg�&�gl�ܛ}
�@ƒ!�������O|>N����ZOD�F{�1������q i�.x$g�a}�+7'T��n�2�jT&v?V�V���ul����͛]����?�~��+�|��s4wBl���"����@1��e�m�3�-��J#�\|�xO�Ii�z�ݿ�A�RtgOჅ o�B�I.�G��ׇ�&�pw{p��Zw��	�kc����C�[}��=�����S�u=�����{V�slCI�aJYD��Qr9D��k����t�1�
�G��h嚑o~��S��/x��AgK�������rG$�v���m�>�uؿ�(��$�{p�XA�e ���>�,];��+ͤέ�������	oG�E��>��l�H���@+�f&��`��tHv,Cv�Ek=릶op~�-�VѾ�Ru��iu�����~�d�$���Ɩ���ʞ��~�G�q�&U(��n�����I��	�h�7!]�S�������n���*��fem���[�u�%�(�b8�����zg1ac�{w���`�I���9�hIkH����\9��S��:����?�&fs�nH]�Xc�]���?&�������l�Lb6�{��f�Q �����%����5�̙ #�a ��6�!������*��cr!>k��~�j�vM%���sk�B�+Q�u#? �O�E�q7�'-�j��[�G��ۛr��1�
����z`O�v�O���M���V *Vѱ}S*	�,a�#XX��u�1�,HB'��X�~6����>��R�9[ۮ�-�Ȫ2y�6ñ`�>"9:��F�K @����a�T��a	z ��-� =��I,�D�Gml�� R![3�yE�,7V'@��Hv�KT�@�g�(���8�qC�j�����8�����a���ݐ��g��` ����=�4תhi����Lu#��I��T?8�N���RR��
����X[�늊�p��$��s�a(+OR�3������0�#�[��s>q�u�N�����@� ��0w���\O!��Z��jT���~Ìz��Qp�X^�@���r�����u���#=N��6���b��������^��~���.wwwdN��]e#�\翯��3O�}�[�#�vsrrH�,��V��_d&�^~H]B��ȅ尀[�ޭ��`E�eGnS�����}J1�8�R�� 6�v��uuڜ?^� oT���>��)�/Ϻ��^������ݯ��
�pMs�>�YI&q�i��zf��;�"��ퟪG}}����)�A�\��?�_`�SU������S-rl�	eW��4=7�l�MY����72a�%���e�^B}I�z��V]]i�|Q�ι8k��΃fE�<�B��l����s��߱�K�Ijtzr�]wT<�רx2�v�f=x��z�]}��G�>s���Y�	q`Uͱ�B5�O2�e}O2|@�t�P��H�
y���M��5��F ����W���6��'�7 �$ wUR$��i�۾��3#�Ę�<���m�^�tpX���0,<Q1��.;�Ǳ��4: >Xv�E�H�]9R�,/���s	ْa�N��S�D��Q���h	wŨ�X� v{hJ��ga�xP����
.
<~��auۖ?G@?��K�i,��`���3���ʘ�ɡL������E�53k���@����� l�M��sX:җR�+!Jֶ`�a��ں��ݶEq�Lh!�5�@eZ��y�s�?������3w��Ec6�O^���#�k�!;U�'����t·��0[=�af���VP�>��ϧgp��\�gU�`o:��r,<ƚ!p�����V�V� ���-�>,i����L���*萒3\}ժUa��ݟRΞ�4M�t���nn���A����X� EdN�=�Zձ��;�d�[��"E�2W|�"�_�ڃ��7��3�B;�v��V$���2�g�0��U|2Fx��<`Eb�R8d(VR�\wzgn�޸R{EEE�3�9���ت�.�XRoo�C�����X>B�ta�H0̫J؁8�e��,�ׯ֠��/g���`z��� o%�q��[>����+(%}pݳm�X*|I�?秗�� |㶥�z��#p�X��/{ �s�`�B�P:�0[�V����((�vk�qJي&��c���?O̴����İ���A�)��1��[o)^*}����驍�F
�熁d���_�򌑂cYw4�3�߫�^���R��;0�f'm�-ð�(H[<k��7$Kig&ݚ����+VbM�P��֙�"��x�ǫ�E��p�	�Z�9fd%�`�Y��l��@�W`4�qSS������K����CJ6ݓQ��z������3�N�ݽWz"'V{c��@���S�ӻqq�}(҃}�����X�'�\��a'N��r���OL�4pkȯL����,{3BAf�lT|����7q�8{Hw�br���B��O�1I�B�rq|t{��ͫ�����[�>�ڊ�
�a��p/��>�/F�&1�j��o�4A��7��_bui�\������x̻mL� �Xp�����ɟ�\$6�HI��'&<�H)m�{6�5�d�����*�"�y��j.�]閕E�:�/^���NFõ���஺��1d�%��O�s�*�F�����[�b�TG��:;њ[$D$�`ɍY��M>ǭ�C'{����,���b��[��R��?�5��AE��q�M$J/�)�⩩�ɮ�(�;6'��K�c`ا�y��}���U'>������D���肬��J;����Gs���)`V{r8� �AE;��`�d�7��"�[>y3af-ƊR�BW��g��}�r|#G�4}�S�mY]�1�� 'B"35k�0"������h��#G4�1O�*��mT|���Q����)�\��/��D8	�:�I|�fR�7�������$[�����Xb�z_������'�r��q�/r,�����OÑc?��Qי���U���R�4gr��G����D+M�<|L�G֎�����|�k��u_&��6a,��f��tyhF�^ئ��-V$᫴A��2��k�EX�ǫ ˃E �x1�؞T�=�d���w�;t�T��khb��������e`�J���5qyXy�ׯW�ə�> ��ز6v�C����&$�9b�l�1ep���Y��s��� 64����QW�c�%��\���L��j'��{�E0�G��h�PY%)fy�?7 -�L��$$ۍM�/n�`|/���b\��9x�qT��︒^+i)1��� ��寧��q�PD�`>��s��o��uv3��Z8���$!�,'����VF\�$������f:0H��� �M6������]�Ru�g@�����0�����%�y��FDDL&�N˦�p� ��2�����.�� ��	��8���N�3Ǎ�mL��1�($��$;� p�r�}���$�4�*�����b��`�)���) 5$j�A�A1���7p?���$_ct�Iʼ���_���&|�1(�z��}�}j�J�嫈?mtq��m߼|�����Flz	�X߳N�<דpT��N����;��lߺu)�DD,R��^�g���D΃�(>�E�𭐦�j^J8ؿ9�|7�O�'���8��H:@D�6�jgE��`�_�Xb,p<���w?�3���~��~�cRJ^��'N��XrH����[44Nݓ)<."���AV}�ƞ�+�]����?v�'t�JE���I`���l�J!�Sp��h���<f�#>|����s�Pd��A(9a�x>�(t�PAK$6
v���^�|c6>Q�n�����0snyqV������KX�O ���̤�Gb�\�`8����1}K�00ȨCZ쨬���HI��ʅp��'������:��3;�u��UUJ}F������Ea�D#�>�G��N..8�n>]��aqiVqq�>�'�q$?>��Q~ե�9�J������ڇ��@-���JI�`�ZWy�ӯ�⭩���h�w-�>�ѱk;J9�m����@�QY���¢Nۋ8n�������nә�J�q���9�W���(���M��.��U`)��Ҏ58�aJp-	S� 8KU=���������g�U��G���~��''\3Μ����Kx7�|�
Wva�S�<��B�z��p��E�V��;w0�=��t� �֙��@�ƑaƵ�=�C9d��.Nȓ��`��Y$�T��:�����E%eP,�׾���)n�}H2"���TYk:�N���%�Q4��n:�ࠎP�QX�i`�H��ppq� �f������=(
��Qd���&�Iq<��;=}>������  ��6��FC�ٟ�B�>oo�Bug���y��m1L&�)�"@��~���~~����DIT�.�ٕ�|/p��Ī&#`TLbPܠeE|��Y%��sG@��MvD��|����z��f��k�$[�̰�ޅ��UD �`�4� ��fq�*� ^e$\� \���˴r ��e@�[���mֿLġ�ɲ�|�C�̲����X�0���*���:N:>��Y�IW�������W�]Vf tN��G�k�뙌rlc��3�k�Bb��ʧ�_�z��P�2��iy�����	''��ER5�7�"�,pȵ��sk��c���s�I&�����Sˮ��w}H
8�������������)o#�	�iO�������_,��E�߭�zw{��[���O�Q����R�f:�q��H�@�I�[D�\�]�w�7��i��k�u�|�ׄ}E��Nc^�9�Ѯ�1���`���V�>���c��#�9?r�4�xz�������ή1��e} 6XV��	�#Va��`��� �J �/ ��Ƽ�;����yȑsR[�ۓp���"�,x4��!����dm�ٳ����t��Qr��(1|�'؆	�6ؿ��ش�h���=�#�(�L ~��\SÁ4�2^������� W}�;l�"v�H\�`%
�2�a~6H!�;�ٜyʅ�[�6�V���
��^�ظ#Z"��^^�!E���v��H�A�1L�\M�;?v9����{��ar�a'���焽���\*#��;�d��4�S��_���CCn�{���`[($c�� ��k�]���p/���ׯ㳷�&xB8��7%���P������ɥ%	��OY�r�)g���`��:ߑu�O	j�>�'''u�m��6<)����?���l⬓SYm�L����,�0�I�H�ryp��B�BN��e0v�$���5@`v�aɦ{��/��w]3���8���� J�?���t�;���㲈Uj ��R:��u�S-��+�����/��NI@^��Ȕ��/vg��/�S��ؓ�e�Vw��֒л�zOFI$�[]r����1�Vdu�)�����ս����	(±��fb>)_�}Ѓ��ޛ�s�}��*�I)�d()*�A��TH�d�P2ː�ӫ�2%EiN$�1D�d(S2� e�Td&�e����W�܏���������p]��kx��Z{�A9^�e��2�����x��uUpD{g�[l��,��2�g�<y;a�s�ў���Pe]���]�|a>�bn/�d�B���9^M&��=n{��l��6�������%�S���~��˻�.�c��*j�ˣO1-AE`��<
�u�c�c��AgW{�P�7�YAu�0����
��:��͍�#�"v[�J\��kH�f���2���l�f�[qջF-`SO}�&������>��g.� 4��9�K�� #o�C�M 9C~����q��#_D���<��Q��"8��:~Gy8
 �9|�y=�*�CQrt�\)M�)]�~ȷ7i�\��	[W�/7o�cs��T��9O�Rc�u"�"�Ї���s��#C���I=R!ˋ?������|i/��#�_]^��5K?2�n4�wIRJ��@���鼊��f$�f[@�ld[q����%��̹؉Rxm0� ����*ܳU&Մw��l��������8�_���R@����솻j0y�r�0���`Sv���
G.���1��-c]<�jL�*�j�Mb<�p/ �8����	���;d��ݰ�  �%r&�c[j� /Nj?$f�?`&(aXsl�Ȣ�l\0C/$.!�F�dm�%{�+��X�6ŋ�L�^B�+��6�Y�;q��$ŅNܟ���*l��}u���/��U1>B��g8�w�h�,��LO�+,�=�[Uq?�$dF�N��ͩ7A��`���ǞlC�7�XΓh~wsm�r�	���A�\::H� x*��$�ZY�z�n�X����Va*�-���k�3 v�������Ǧ���\Cq��'e���,A��L�^�(� w�#�K�b���x�}T��?cg��V����s��#uC
ˉuuz@��#��^¨A
/�t�?���${X�W�n���V`�׎�&��ƾ|��t3�f<ݧ�:�g#^�>g�
�����oC�o��__��l�&�����l�6AR��-�0n>��O/���j[<`��	*�Ǜ}p>X\���^�(�gcɤ����J�T�	6!i<�F�q-�`a>�B��[d��LOݐˍ?���M;"��}�J't���j$jt���������P�@�v�7��u��Ⳉ��z`g d����3�H�d���uCzz�J�˱��?���A�*��nڴ	���#�i�[r~�,�?� ������emb�z�lP�o �>�4jD*
`�]H#䭿�6�$`�R��h��:���!k"������W*�Y�h�㌝�6^��h#�}���y��A�37� ������&�}�t9s�^�~k���\Z5�n�%��m�6�f�@I��yV�l�y�e��3�ϱ��BΡ�<�}�iWf���F4?�1c��7��.�O��\@����K������;�0qxء���ߊ߉i#^\@_�w8INYL
�J����+���	��{�g�ݥ��6<{V��*Ss�������rI���m��c!ۻ��ѾFb�o�C �_�a^�Q�Eړ�ӂf�P�=��`^5�ޞ�-��k���3L?Z����9OH���8��h�	!bݾ�F�B�����7�QX3r��m��;���n�Ѣ/q [K��G�-׾�Wk�|��������� ui0g�����I�J������6CxōZ����qTvKP���C촋
���/.V;ʶ��%b���mHH�[�ı[�0_y���S�>vYP}BB⎯�<�;�6�8a7]\��UQvͧ�q��h�$�D��$�^��\�_�B~�|���:����v�\�����V���qZ�o��h��j�t��X���Kz�r?�2�V@�F���G#�a�ծ�w����J�}V�j��чuY�^�.�#t3q�G�5r�u�7}�����Pl��37�X����Ѱ���l[{@�X1(o^.������<�r�
G[��cο鄹b�o���S߸VdC�����Q���⍷ߏ������g5�����%�V��=��=�Pc$�ddƨ_�m�˾�f���I4Z<Mmu�	ZRJ��٭1��v�������+;�-���/��rzwt�����7��w����S��L�}�(�F����|��[� ���>�=j�=�>.�@�o�/!��ؘ%�܆�&�Ts��ֲ���]���ߚJ���TI��y`��n	'6��x
 ���Q�L�ٳ����O�e���jkk�������[�c�a����_.�:I��J���Q���i�Z���KĄ����� �v���x<�����I��c�4|,�V��~R�G� �y��w~~�}�"���95y,��șY��)�8+"L�/��06����zu�����\SkHk�54H�n`�t�+v���S�J�S�����8��wR��[�D_�N��X� '����!ɷ.qV�i�: ������{�P�����U��s"ה��1��S��.g�a�}�؇��1�������M�`cݟ��7�����}�Ǿ��J\z��iÔ�Y'���[�&��TD`������7���o����CFh��pu�#��a^����s۷�3�U�Va�.66��[3Ը�˗B�����ԇK5���!��x��6j,b�4������y��y�
^RJ�����p���	Me�չ�`�xa�ٽ� %<��t�1m��k�'*'�vX���u0XZvO�NO{��=;㊭S4�I 2vv�d>�FG!��SЋ�'��]-��*�H��`�T�m��|/8��]Lxz���g�P���y������EJ�r�Fg¶�����W��Wm�(�qqg���]��^��m';#���!W�����47���́��c�OާO�l��r@��I����tE\��|E�DN���`\�K9��ܥ���@�f}�Jn�P��}��Ny�C�@�$�a�&�c+b�G��Ɂ�E��� ��o�B�s�d�m�����p����Y=��j��	Q#G�T�ݲ u4�7��| �Ӎ�׳�3��cw��쟙�Wq�h�� _qz���c���c�����z�
Wo�d*�Xpv�
�^�G��E��M�N�}�ä���Ub}��77o~�v�P��,�턹��v̴sw�6��-{�B2\�H�o,e�!�s�4Sp��ɱ���-�+ ���XЧ�!�����L}m4������!1i�n�(�J���Ǉf
�� Sx�6�����TFV�a�����C�Ş��lͦ���:�����I��QѬ��/>yg��=�ۨ��=āM^�Sb�5C(5	w0qP�GuC��s�S��N�:���ϱ�{4##��ƁK�T�I�uڸ�8�zId�===�%Mǚ��@�lW�_����Z�s&������~%%�'\a/�`3�2M6��O�G<a�}˖-�A^��[��FB�-��]�a ;� %�?�l"����`�\�\���^�	��鶦�є� ����\ӽ�[��HO���7��1���J3CJ X�Nn�z�S�ӨW��SEsT'�~����]�;s������{���V�rD���0�]�x&gI���[.�`bb7�����x�������%�y�6ɠ)�*:Q� ¢�<�A��҂�5K��t��t-̭Ou �R�?��P^p�kRI�{��b~�A.�u�#SI��_��{�Q���v��c�{0��7IH@��J�#����qϋz����ё#m5���ț���8*�/�O�7R=��J���U�S�S�fF䈗��b�{�Lv�%|�2�*�;���C��|�XqQ�jU�1	i��4�tg��3�J32��
S&m�!���������~��aeg�ZZ�9M��=%J~L��6��.�|����K��Z��SI*�,rrǌ�������Ι���K ���!J����lQՄ�=����'�?gF���>�"~/��h]]�����Ї)��f��FMs�XL�D6.���䠜����نk��=tF0.�q�[)���3������fk�LufR;�f�+{��,./�iU�m�ZZ��&{*���*�g�q�O_X���!b��Du����������Sl��M+u�5KZV�@���ݲ���!�P��2n�6WG�'�Ѡ��UTT��u��І�H��'qq@}w�ޛ?��0ܹ�t;�u�>+b]U}��Y�`���678cB<w~���Lh��Fƹ�l��ԸC��7�p�>����p�1jll$�1D�x����K܋ ��C����8-�C�U����������|�U�+�Y�e��4	0��epZeM`l`b�����k!����X�O���ߊo�r9VaD2�-//'�a���&`!���o������kP��ݓ)��A��ޜ�����~mc)�)P�B�u �O*�n�MR��˫��FD
mȵ����UUUx�4(��-����NBn��2��\|��ʁ|'��F��'�R,B�=��>���C�7����KƤ�?�5\[�-l��Q�I��J�\��񻀠 �:Qg�/�x�2�������@K$�
.�F�&絍��:�}�J޾�|������*�s��f�Kb�O��@���V้�������K9dV��+��K����@��`3&` tw^3d��^�u��Vp� ����e&D�Lz��t���%��GFhm�E椊1�n��^ƅ��k�h<o Yy8��w�?v��"	O3�
<��۵�7 ��G��Zp(��Vi������ǎk-��l¶Tħƀx���Y�o���i�]]�͏���*���!����ߨ\Qp��?0�Q�� Zb<�7�k��k�gx<;��ٕ��+�%ﭰuv^��Q�i���gۓnYk�s�s[��3�-��1�)U��u�6��(���� `�t�fmmU��0fy.����Ĥ$$��-7KMRW,�������(�ѕ�{����+��8Y��*�oE�:�Z�ׯ#�l/\X��6�J&.�s��,5 V
��7�����1��t9�	S����W'4��ׇ��]jB��/%�+3���!�ѥ��Ee�8`Yiv�!�0���a_��`�����\ ���n��:�3�U�ir
�'��Jo�A��%dP;Ƞf��?U��$Uw�o����F�v�ăi t������;W��0�l�$��*��MME�_;f��_�E�� �g�+n�Z2vn�<0�s�0��s�v����ϙ��ұ�]�J���X<��xt�����8?�C�$�Y:b;�	ۯzx���,�����B��m#�����bH�h@�,5���ZCK2��ƒ��e�A�s.� ���sK;I�*�-j�<a��%J�d�}�����v�� � ���'��99�%9�4�]Y��r�n�6@��e�:�$�-�,$$����,}����ʉ�4��%��O�c{_g���y0n/�=��������\��`���JB�y��Ǖf��o��3�[��}�|����XH'�J8�na�O�ã�@Ǻ��h>��5a<2

�غ�Lr�&���qugv����	R�~!�w* ����	,"/RS���� =��"�(���1<���ф^#��wlU�����	E���2WG�;�O6\���e1
�Mo+'M�p-�0cͳ  :�Z���>���һ���uķ��� J�ӧ!�Y
IIM��*6�_�{�(N�"!��Z�	�!�,��|ym'�1x/�[�1�V���K�a�F2;� u�p�
H5w�27:�`��,����Y����B��V��,E�ƕ��s����2�~��$FO�^--/I���U/��nӓ�����z��,$e02����g� x�H������_<�`�+H9"7��$Kq#��EG@��xW�  ��U����+����[��?�˗~����G��%du�����C��cc���~J
G����^m߁���&���,��-���V<j���}�>/��I�w��T��5N����+�x }iT�/��
F�%�`�Je�	cx�i��J[[O��l	�c9�t-�/���vᎪ��K`Q��uR����	�|+/?jzc�&�i�)��@��\����#~-��~�é�)gH��,����(����e�J �%��<LO�8q��7Sģ���X�� sU�r UW���F��)�N�������iG9�we��� �� n�Eg���j�����夑�\����=�N{g��q�
����;� ������=H{���#a�����}���P�5���D��1:���iU����H�r�ӿ�,x� 2oU�g>�J�T<I/�o��|��Y`�@V�Z>dxg�o!E�\�g�����%�'�7��pu���]�v�r,2� �t�"���k�"	�6|�����\@�ae&��<"��O!�Ӫy~�����j�&����Aꡟ�.띿���@KK�v�����#�'�<�-n�wl����q�0H�8�"+��_�xC'�6 �E�#��2�v9E�� �+E �?�>�j���������¬���Wo�n�G/�����}V�,e��	�_Gw�cox�|Y	^m���;���3�rEfkXY���KոnY�e�x���K'�b��4+^��(n 8�հP�q�9Q�"Ľ��Q$䬇��q�y���`3I>�3 O���p8]96&G{MGB��E���!�C�`��J�K�>`�ԺV����H��n��/�BzO;�5�3�(��c`�aR6�vF�G�Ed7��NC�$�[�
���
����\��[Vv�$�~��x�߬���&�'��h1��MP�/6F���� �j�)7
���v��("�(�Q��7[���Ѓ�Uq�]���f���J� �#/ �� qE��?���5
/c�+>Azx�3�+2Gy�NxD#=��OPA�;
�I��7�S��d��k���c-mF�yo��퀡Ĭ�CROa�+<��BNF�m���&�o���'���D�v�����(��4's�O�L��`\\̿����~�q�kQb��?{/�&b�1$U�����.��"�k��^��A�#�+��`3qjο��|jlLMM�xjd-x ��9�5��Hv��Z��E����Me�]38Jf�"��L)"�_�1���%�+4T;���3c�3�u�����,--+͜}���!���NFA,C����@�I�p<pr:I�������yy5.�J
�����oQ�'�o0�.Ƒ���c�U[���dh}�x寅�u���7�Ga��4�K8ede����@&� *\"T!l�$��v�0�Ҋ)?��fUVhG�%(��A:�#��K@rC �!Ti����'f��X�b�-$�h�g�.#���?�x���{�ǝ���1E�X�֢]�v=h�L&��=�j��� ���L�Ϩ�V�ل�ᕤ���0rRi�v��J�������Ԇ�H�!�q�X�3�k�c��	��,���[�J4)��[�1+ވE�T�����d-�O�������Do�k�<N�A
{�(p? �f�rU��p���So_��5�+)��K�s�%M�m$��ؚ��D�*փs�E����'��*�1qq�.���X�`�<blĲ$?����ׯ�w�f?�&E�ܫY����"�G��⻑G`�c0�+^Z���y+��@�ܧ����:�I����h\>S;�*�X$����}�1=�Ar�:�����$Q�����?M������{{����JLI����`n��脖XDJrx����om�
�T�E��c'�=���b�������z�R5�Q"�S�`�U�l��ռ3X��6���:`�~M>�n����0��Dg���M`��''���p7�|�[	�s>����m��"�K�@4a ��g}�o����L1UUU�Bۿ!p��U!�
�WCvg,!d,^���$��U�5��e}L�,'�;I1JR�L�(�k�*ͮ��]�sy�����/**J��kt��$�!>����<`�1f�:Y�EtD�`�aˍb5~!!:y�b�I��k�u��1��s61I��Ŵ Ҙf,�n��/I�z�k�Aas�%��F4����v�B_��*�_�>�̄4�15��+��������@�k��ބq%���?1�O�����	+;��ފ����}*b����ԃPn(!LT1V�3����ݖ�q��.Lu��$/���"��.KY�=(Cs�F�8���Z�MS!�O	��b��Ak���v|�?��(I�j#	�"q6��`�\��`	���������B.���� ���Gd�#�W��FRg�bjE+%���W=�90�(�,7�/��8�-!�Bc�%gf�����c�98Ԩ�!+�V�%;�y�����!���� ��A�c���e1�M�K-��<ʇb���$�� � >��:P:욕�����m�DYwl��T���"q=�ɠJ����0DEX�8�\F�/��&j� j��z���w�Զ
SH����VA�$%[,��72R�A�6#-'GZ@�$V�^��>"%6n$.Y�CT��1Sݞ��B^����Aa�E��dX5cU�3�\�2=+K@JJ���U#�B��P�䙳������Y�7��c�.\h�m���"M��xK=�,��PN�/;\1bymX�9J9C��UN��b���lJ�o�
�?f�=Hl8��J�~KW�Q�\�c�p)
a��l��$�zP����6%�؄# ������BP@{i���8���(����6؀��BP�NW줥����ߣc�$�L�%��Ҳ�׊�HKۙ�9Î�C�Ha��%0�f�����~����FOlU�7(4G��S_��"N���V�"8h�H���Li��w'�8v�ZdB/�����D�����A���}� �D�Mi�cj�奄/)�ȹ��*�C�wᕗ��|�p�fS�v!γ�/pF|CEܳ�����g��">�=vz�CǼ7�ͳ��W��k%.� �܀D�!l�H�s������tv��Oy%E��Q��g��5$5��>���d�(sQ��-�L��/Yx�d�$J��G��"-mR��ٺ"�V���\���vzu�lF�t��L�Dp�1�#tn�"g\X7"�2�F�v��]�j%á2��X��z��>@Fgt��"T�� �X��ǀ�zV.���){	�r�\!,��u_{N���:"���J<&��A�� ���W��F��҂���]�3oz�O(K�m��$��Ux7��<�*4�T���ÌΦ��?~�xmb[۠ta�]��S��v�~	�38��N ���5���c��![�8�Z�F{�N�ʝ|��JJR�f�����%��®Y�]<��Ț;K1D��a�.пjHЕe��]���d�Eh�.3�c����A��Eq�B�*CȈ_JKKH�Z^�	������|�qa�ǝ�G�g�������/��kSI�� O���ZlE����:���c�� +��ۀ8���}6�2�4��x?f@٠׽�]�ꩫ�c���0hç�%,�)M�,B
ڑ<��6y�J�V�a�0Se�+ h�K?Q���ܖ�34��}����~��i���J�C�	��ڃ��TH���(�4d���Q$sI�{���h�ir��L�!+YE�>�q������2�Y?�����%d2��*3I\�Ɣ66�0"�v�k>���K ��Ҹ+?�_��7��F,��M�HI����u�إx@��6�JA;�|�,FAQ�d�ü�]�ͫ�s<{e~�~����k���fiz����9|;[���I�)7Bn	�N����)�R�D��ɇ�(C}����~O�K>ŚP*�Á��{�G�*I]r03�aD��X�k��t�:��A����{�$�����|�^�,Dܢ����gx=����/�I9�u�wE�T��N�p���i��VuJB�$��.=3sUGGD��L�&�����l��H�|������O��_��yvʰ���J�>���xi���T�!)��,��XЏqKO�)��#���F*5���ʿ�l)�5kc�U���8�[���I#�}�����R:4 ��-r`��(�r���	�-xxϋ(�
�
�����q�؁&�!�o^ņ����,�E��7f�o�:�eu��SSSg�Hd��|i��P��a�G�,�ӌU/4�xg+�z�K��>p�YYS�*<��#�lr�2�6�a�ƤzTK��@L%�ʰ�EԁJc����&F����Ǫ_r�sQ6�3Gh �!��@>^S�a`)��/!�u_��%�(�zz���p�VB������k��#�^ͥ����tk7܂� `I�r=�u�@�9�� ����X��X���Юu�Q��Qr�+J~��R���K����I���"�.h$���a����[�m��&v�=�wMJ�-m6.���9��msl�(4�;�D༘��տ-�Z�¤�s�6O���<.������+��0  3�r��!r�W�ެ�k/@E��5��lu��$F#�~9��tj�tA�_�$c0���`47����'�����>F���^S�"v'Ւ4Y��p��p��'b�w�c�l-hd�"n���P��*fC-�����I#��zf}�4��D}	z�}�Z����^����5!	�_y��am7�y�&m$x\&�>C���.�x�
�+}�t_=vT�����(j�F\\����U�v�~��&���`����� A��H�䏒wC3E_¥�n޵�|U����={�S]JJE�}u��2y]���/���)���w(>�U��|�7ї���X$T��ei���u�? \6���J��]�2=�����ז�7t�?Ej,vN�Ux��V�6f:W\R��)}�p"@|��*��x�6zKav��D!O���T�\"��Z�3s �G;���vh}H����W��+�6�>Pm��1Xd�0�{�����i��%BE�pA�͛K�(��%���p�L��T��aW�S�N�uK�%��XhM�S��7���������'�v��{S��8� �ËY�$�}�X��BH�AZX �1��X<2��������':�'`� 4�4��b��Q�w�)DS�mD��sHs<���C�N��mdc�L2��s��15_��[<�07��Û�l$n/��u�*A�3�����:#�L�jø ��"��P���C|��7&���	�Iϑ��P�%�P�Y�d�s];I���t
pZ�c�5�)���|:�����(17.��ABJ��+J"�is���蘩��o��p�u[a�4�-
)y^;�$Mo���`��!?��:�[�vƘ�A�{���낅��#���Y��L&'�f��jD��}�o+�R��Z�^B����Ρtt`�`� �!ŏzdl7c�=�V���$ƌ0��:�'$:ȕ+":/ꍈ0���]XF%�0�к����K�F�����+��* �m���� ����`�3�Jv..�#"� ;�o?�����2��ڽa}��!�V�Y��o�򁖱^�h.��\<�P�4Ïņt��y6;�YH�U�?������?�0^ty�;
���aEAB0�M��r#iw>,�ה#��6B�cc~ˉ{�<�t�聘�`�͡��'p�K?,�6���"M�0i�{	Ћ6�$���g��Szz��Et��SD?Ⱥ���m�T��ǌ5�}273ɘ��Nx�o��%I�YK:m7�G��K�F�<��C���	*�8v�#B�y򜓓�g��g6&8 .�WD�%���uU�%�-��<s���\ޝ�H�g̑���db�A8�S�^EX�0�я�����C�������[!e�T�Y~�ۼ,��%��̆6��b�����}�Er&���3\�v&^B�˸�����#�>��ȟ��3=�	��mz�K�y-w���؃�cCH�A�*@2�_q�
���9� m�����O\��<q"�-�5���^@Y?˾���PﮉTOi~���n��a�ݑ�ѵj�)(�S�h�p#M������wY	&���̮5 �''��eK6�c��gom��T,K��i&���0p��Wq����`�v��s�7�-ix���l����ZG����7U�oZ�6�c��G@S����ү� ��!���A�]%X��x|ͻ�C=\����nf��U��{d��Y��ↇ�i,tw��2�|�g��.�3]��M��#s>@�4�@tI*���kˢ9�����OZdv�}���W�7���:u����� @!	q�� ���^e���d$��Ѫ@RX��&���f)Ms�����vP��_�%AN�r���0��ԭV��R����8s�M��)H�0|���'���Y�d�0�wY��,2�w�@L�9�|�?�j/�d[���"!���-fv����v�NNU$�̳���
h��J�|�\�ͅ@���:�{��?u�0�*A���_ =﬊�st<1"�#]��3䓇��Ӡ���Y��]���d����@��~��`��RAe���״<���5�I\�5��OK�FE��G̡����Ō��B��q�װB���.#fм�.pwL[pD.���� ��������l.�d�E�"_�)	�5��[���+k�����mAJ���v��@��`h-egG+$29r�o�^R,o�k�q9�&�i����v���\���z�~U�F����1�=_Ԇ�ށ+�P�+�߲�.�7��mP�����,� � AeH?萰g)�� � ��G���W�7޼���dI�2�e��ǚ	'�V�k˳�H�*��7y�lQƣ����ٯ�W-_L^�K����']����,��(C �U�=���-MoY&��x�|�����7Rz��B�£�4�^%t�����u�
�<n!X�My�����5+P%��WAp�v�K�&����iy;TI����͈"3���l7c�	��qm�ᷢ�.�H���ř�� �ɣD\�Z� ��h�s���:��E��@�4":�[��T���W��]����`ZP����;�KD�7碨F�;���bXj'նuDz�N�@8���m0$i~�(5ŗ}��60^v^�ktL��+70u1�[q �$�#J�W�z��2�������k��v�-��z0{0�T��CT�`8d�=��UO;�k���JH�M���R���f��mX��ى>J=~�0�K��g� �>V�_#�Fl�!����g���^�x19�ɰ\OFh�]����˃���e�-x(}���pIʻ�R'�:�{�ڵ�DC��nh���M�6NcU�cs<2��n�Z]C�$b�S!� 0L�7��E�`|.yNo-73�1�5�?�xs>{�L����2�D��J~�;�����:�(O�|�5_�ˠᨣOo�^�l���{�Q�������Q�
����?�Ց�@�^H��xB�BI��@�c���l�90�E�435V��ϳ�������b񕺵��eee�#=�t��{%�\��j��Ǒ����aw��$^=R|�5�3�������EYڄ3�i���{��kz�� ��}����>xq�&y��[�Q���m�\���O��0״�e�����X�ڭ�z��:�d�6 M��1|ÃA�k����-�+�sO;G���<�ٮ0�`�f�t�r�O�]GZ7�EWu�uT�MN��Q��pmQh�-����r����K'��,%R������8L���i��G���\���ϩ�Cμ:V`�@����g��6����xۿY@�"������������^_��5�n�n�}o�V��pw���3aj��Ly� _p05�P���+�2�+ί+�In A�P@Z���,�;L�W�h��x,-7�g��Dg��fɄ�s�i������9����z�{�>׀<ؔ���~RH��Ã%6V4H>��ޫFkw[$$�NyW$�U���SqbqGm�E)�)��u�x	6�ϔ�����T3܀7`��+/�� �]bH���������o~��<��r�)N �ޚ�*��:*���ݒT�V:/C���KՉ�"��OOL|�YJ0Ȉ��|fdn<���R`��q�sA�������+1�N�I�r
(���o����(�X���X�����5�=��S�V�fe��sO@��y�k��m���:����KQ��t4��%S<�����TB�é� �6��lZX���('�Ԝ$S�m�=�������)��L%���L��N�R0-$�3f�QDט�wC�X�=�uX�p���G�i�Ne{F��|>m�9�?X���"b%�C�ש����@�M�����C�_���n��R֜lW2i����P��Ѽ�3#�_��s�R9�r��˯,�J��/ğ�z�c���'Ob�m�6�0��\޴�s��}O�DM�im�%���ڟ�:0O`kR�UKKKڳ��ӡKnM�f�����|!���W�>��3N�S�����A�L�{��' X��W�%�J�����TyMn�n�Vr�Κ�y���٬<ix�9ٝ�����_�'5W�٭$E|'��w|�R|G(�d��.,T��VȮ��@�O&�Ú9n5�����9�fƌ.+&�w,�d�>��%e`ȳ��#}	�V��\9ଂ;��k��d�!�gDg�0�E��F�3���vG���آ�ɫ��)�Ҧ�J_�5nS
��A_��d�r*���ib�6�BI���P�Ӊ�;�"?t�X�/�����&�@��!*�6�ed�9�vZ1u�{���)R��q~�?�#PBjb���Le�'�`2�����ي�]K�>)�Ԕ�%J�{�'��0^��egZ��C0��63|�C0� ����!%מ������L��e�=:�cCJ+g5��^Q쓤�ن�+��}����ր� ��?��0��a�p_�¶��;�7#9�# A�[���N.;7Q�$��h�ck�0��y����k� LK
�����<'_ I�LMMQLL�����rN��3�Q8�`@��Gy�~�	R��N�׮�i0�������F��c�n�5;_�~f��ڒ�زK����9��x+���M����q<����%�S
�U��p�
g]��G��a�	0�+�$ݙ$��9�Mזb��_qP���� -���b��ϓ,�j�x_�X[�:#�-�8/�G*�#�n,�
D��Ӹs�v��>�N@w� F��p���bI�V���@�9_}}=� UUUL<��n�?`7���vT�v��U7DԀ��bMK�n� !�/p�K�K�A�|Q��˗.rBD*��X	q�U	R7�p��ԟ�R?dAH).V�GG`��@FF������M�ì$00�M��5P���.����XV��V�ؐ���|���KOw$�5�Q���AT3O�"��MS��I�J�y�`eaRv���#�?Z?S�>9���Ql�hw�fAշoƨ%H����Q&����������<2��gc��UL q�M�{�.�nF���4ˇy�S���b�ƀᠱ�����F�T\W��JD�.��6;��=j��Aqw�O���cxdDF~$�d>hӐL�Oi��:~�q%����sJ����h1�&D�̳��Nb�}z��L�*;�|˟���畃E�+��3�e�@�If[��ص����`�;���y|���Wr5m\�`�Xn�A5�>��;|�N��r�a	#��5�w
�CC�i��;s`עEѵݷ��67�u/ʒ�!nɤ2NГ�[}�
;T�:"`�v3�G���Aʍ\�em��\��_�EؽG�oۊ����\TDF鄝+�[&��thg��Ss:�p���X$����Z�bn��@�-��j`�����藎�x^��(k�RXH5�?��F�
�b'��BZ�w-%����͙N��@J�	��v��#�C��>�5j&�D|��7�cS0wT�k�>Z��m�΍�R@��O��V@�S��	�3�nӃ�(�K��M!5��1���4c1��U��ϱ�
�ɧ ���H�\3D*��s�58(�y�y`�(,������4XW1�}�����k��E��0-���!�^b�X9�x ��8��I�V[G�I�(��n��..���io�i��M8�S�u�O#�*c=�*{�v#�����LEz&�N���K� kH�Q�Z@  ����֦1�J���*�cl2�-�6���m0e���p$^��m�L����۽�����9~���o�c��q��^��~҂�ر�|���O!��	����R��m�~�H�O�
� ����V���Y�BOJ��xI���nY�� B#\�XHeĘؼ����Z0$��%i��7wp�	��UyEE}��2xrvװ+X
�=��)���!88 4�I��R�t$9`���B�.yz"q�4�`N�99�����%)�+���<�EDs(�'���$����	�S^�+��n����/����u�V{zk �^On��B�,��5����,A�& �@�In5���[��A����b�-Z�'�i� ��n0L�4��,K�&�O��1J.a}l-��� ���p�7��$1X�fb�3t�$>K��i%6����r.ĝ��0�C�U)l�����ǰ���r��'��P���jU�txŒ����WX��=���k/��Z0�'w��^��}��u��K�Q��­�UUÚ��X��`�Q� [�t��(�i���2�:�����x�Ghg�-��*��J��S�	;X����(�K���h\F2�v��N����C�%<V���fz��t�u����+@M �I 8�@�]D�� �IbW��l�_g7�yiz�q�#�YDV��#[�M�6��"[E��v�<�z0�F	�|.2�->�&%H5d@��� ~����e)8�=pۅ�8��QX����C�Z��F}u�����`��U���"[GGhF���I ���m�ap)ؠ�y�Y��;&HEe����im��tm���fh��K�0�$Q�\��)�kk1�O�����|��ȣs֩m����ײ����0~���CnJ��6R�o�]x� +������s_��N� %w�c1�@�@7�krp������N|N`"f��4_��FFkw��%,�W4666�j�VZ�e����L��jjj0>�R$ӵ[���ƺ�	f�������L��aI8x9{�!�<��!;;{� ����lX@�?:B��ĕ���l:�h �al���o��iM� G��k� ���N��	�&�2� ������kK�7�F�s�~񨓫Ղ]�SS����l������g� ��I�r(&+�e\��g���6.���qYG k����f����Q�~Eep�-n���v��"﨤���� �x Xw;}�*��״�5 �L9	Ɩ��4۷o�o�ˣ@o`d~�
�i��M�s���V[��U[����s��|Q�0��)OeMx���`��YRm7k�bᴚ����d���#��\\Vb�5@\LI!
�f�N?��n�.M7'�D��6Yixd.��]~_`k[Q�� ���o��;"œ��㮸=�|*y4�2��%@aI����d����X�hII	���Y���&6�| �����8�YЫ&�X�����!.�c��uI����b0�CA�C��ݭ˴Ɉ3T]��q~><:s��[.�X�E��Tۡ��� n�QCcNn�A�>��Na�p�`�-���0H-�	��ik �����r
��Y��;�����L����,A�,��^��bhl��ɚ���4�um�Pk�m3�qۃp���Us���tɗ�s�h����WxJ�&Wn�:E^��Ȝ�p�x1Rܦ��o+=)���~Po��F�,�x���ek��s�um!¶Q�]1iu�A^����IW��g�b�� 3��{��Vy2�ě��3�=%܃|���x;r�|�ƒZ�2dԂ�<p|�Ycc��ў���N䀄4ϡ��!�;�v�ח,�No�����*�y%�]�F,���dZ��oҏP��
�|L�d�R�kJ��K>�=�.�J0�`
;���:KP������/����R'ON�%U$�,�Ƀ<�>|�羒>O�¤�6���`#7;��OE�>�t�L�aC�f�k���۾}�<��t��0��o���qIRh��Pk����gJ|Ѷ���X����͓73��m��g���H��*:R��fvML�z:��S^ML�Hj@]��p��L�o�C[=a�d�����l�����4�=�ZSx�_ؕJr;���*2�лm?�Ǌl<��u^���)7���t��=ήT�)�G�c��^��"h�{�e����q��(��gd)��;�pH;�O����/�ݔFO�y�DNeǧ�O$�a��}}�������CEU��3&o�z*�'���D��]١r�Ԃ��Ɇ�5xJ�Dg�/��?�4��h�`���;�"�_�z��/y������I������ǧg��<⾗���8~��v��K�\S
�LL���?.	��[xJR��j춊�;����g7K���vM��'�>��G���02��I�sX�������ڶ�����j�쪭q��rg��gA��+����~��/���������_����~��/����=������l7ɝ;��;fU�|����϶VVW�l޼����qI(�ɾ}V_^���}��Ea��Q�%>��5����2Z�'�ɓ��2^;ILB"Ⱥ�U�%N��������/�	y������;�����J��?�&$$�%}���yޕ=�&�wND(�����y�NMz���w�TjUlEGbU��;w�5�����VY�?8�][T�fi���!rBG[{�����	����KrJ}��6M��#�o�&ZXYM6�	D&�L߲�|�*)k��Ԫ�:3� �32S1�mhzj"��m5�eCCC�<}����vw������_>~u������z�lߪUF5qZL��7��?�)�V�������w�9Rك��?&�+�/`)aF��z��F.�*I��ǿt�Z�&��1�������2:.�+g:�d�ue���
i[C~Of�]��j�MU����v�~v�lzs�2�I�������|~�����-0�c��&e�u^X���V=|�0�(z��<��4O��秕��\���f������'�~	+�CC��P��.�ُ�?���=k��{ā���g����*�q��»5OcW������O�c�ɻ���p9�dn%R[W�WSS�������4-�1iTPD8
�F�9h��wL���\~mAJ��S�6E�EBB>B�ηn���c	,���������1�K���2�d�Ǐ*�ϟ/����	4
R�uu��%{�.�{�ͩ$��d�lF����o4�&���%,��=:��JC�qeZ�gwJ�����w7�ǿG��g}u_�WTo��;�x�����ݩ�w��.�p=ee���Φ�o���ץ��X�M��f}�[6���.������=�my��i�^�(����^K����e��Z��J���ߟ��D��h�ΝxE3��^�����}L����%%mm���)����P�Sެ��km%��?x77ˈ��X�E��"Rh��,`�;+v(���w�o���~Ѹ�_����e�������l�^t����NW��ҲKw]���\u.b�N�C�@��4.�nV�c]��z����sZ�ͭ���q��^zo���[~\x<>һ
�~1Z�PL�֍G5X_l�4��R3����>p���; ���v�+M�A�Yn��
se.����p����r�m}��a~�#�6Ed�Ͼ�<��@uȧٜ�Ά�̷�3�}N9�9Y�w��5"d�i���W�� !!��'z�_F��g��O��ߟ�Hw��xW�F�4BA�W\o!a�f��.4}`���}��닌S�jE����rN�յ�����U��{�W�^�Q�֣vc���؋��we�M��8Q��p�ъ3�=�yg�}������v����F��,@2���?;���c��G���\�F�\~��w~��mO;v;�,��}�z������,��s��˷�:�.�w��5f:�(�+�LJ�}����d��5B�N*jxioT���S�gA��r���Ϧ��dn���֜|�x����Q~/��r����ao��� �
).��V۳���-���یT^��Yj�<��s*�p���XG�]��W.�u�����.�����[Ѭ�[qg���¶Q��*����U_?֨z�e���U���u?��������5�R���e�u6\��J̓�'�ȥK&�bn��*�u~˯cLJB7�=��%^/���pP�G�c�]�;������6@ǲc��95yH��2�p�Y��nݒ�|�;H?���[f�>���}ϱoww�ד�����+���9�����^���ʵ�������l �e�b�!^U��w�Z�V��͵�*3�S�*.e��/���:��Ұ��^�$}�Q�뺩&��e.��r�=�>X`�rey��D�,��'��<�z����n�r��?����Wj�����n߰qR<I�CEH[*+ɸ3J%�(�J��]��)�̌%!��Q�[��##{��=|��������|��u��8��Z����W��?�1?�z�j't���;ĸ��(5r��7IURy˞K�F^�ud �������ZWW�Iw 1�+@Wh�[�S�=s2W>
�B_Z�Z�C�51~�:������z㴴(j�����uU��&�.��o�|^C���9u���)����+_�-��
���S�L�V��X�nU��dґoq�Ǜ�IoY8���՗cB���	�Y&G��Q�̍�A��k��z`1�,S&3՘2?Zd#�'���A:���Pj��ߟo}>Pcv5�;+a�ǔ�'X(���kW������o�	gϜY�I���m_�3g^ز���߾�C��^����͛'e��ͫ����D\�?Emw��|�<5Y���%�~��W��y`�-P�t|���{�i5'���yO7@EY�t��)�UY�			��'�kfϞl�XR�* �`�_Q Pg�]����~5���<��_ ^� �T�|�[5��(c��WDͮL5�2ǫ��Ԝ6C����U9	���p&G����]'x~�����o%�Q�* �_��'�IG^�?�x��+�q!�3�-�ͥ�cc�Z����Uk6�_��WUf�� ��z�4 �Й,� �.��+�V�����}g���w��I�U��T]��>c����6�:ݿn����R���D�f�6I���/���!+�F��������IX�ۘ�&I�S�����I��\��[*��c����@�p�2�p��D�����i�ŧ��툩f;�-���i�w�Yx�~L��ے�D�F��1qq^����K�l���Z'�M�c�ކ���?0Щ_p�l�}j.;QNL�	;���)T{���o��iڠ#&*�	$F����m�� ���A)ɬ�~����\_�S���5�?����̙\:Ueg:Sf�c;�֨�7����7o��R��T����ɏ`����%Y7V� [f�����_�\;z:LV���ϟG)8����jsc���괌�vx��vL������v�lg"N�������y�H��ᬹ�ii�?�xjj[����4�s�֭�Q��{)&��2`�@nQ�S�?�Fcϙ�Mw��o�¶��>�����F�LF���y�-N�hP�Q�p�=Ϥ�a*��6Z���"�=?������i��,jq��W��q@���Z��坖Y%�7:::�%��@�rɀ�IIyP�7a����՘�kHM�ht���yf9̽=�z=%�͕e��kF�M�~>ih������?�nr�FH��Z����h���H�X�#x�zia�C�iV�~�������F�A�x|�+ �t���L�_�R�޻�ϪQ��/@tS��� i?E����)�bov:��.0z�V��
�/w�g��t�wZ�j�cv��\Q�|�e���H�����NEfU�^+�l���9�z�Cs5��K�����@`@��8�Z��ʤW��8����iVS�vJph5���Ϸ�Ϫ���J�x�����y�ݝ��$�szUc�_��SM8�������}ҋ�ʒ����Wiii�b7<Rx'��
�{��B��ӯ�rvЇ2c27��hff�/���w�ځ�<��6���w�kk�=r���	�=��wY�&����Brx�
Yx� j��x�Ƨ@4���	�	�P<[��✨�x��k� ���OX$��/��*2LΪ�ZY�7ݭO؅�!���2�����;=�ё�I�4-�1ABt��Bx�ן�Zy��F�Io^~�칡t�n!�o|N�$Z:�ٷ�)i���T������@�?f/Β9��<��������}_�6�/��	� ����7XQOO���+ �_�z��� �5��V""FC�>+kuc�Iecc�Z���L��t ��
�j�<Pվh�`W6۩&���Y��D��YJP=4�����I���_'Cr��U�޽�.kp-|?�}]
��6�;#��ԡ�L3_�x�"�1��7�������U������T����1}�I�Y�|��!:���@������������z+#"�|9D����k����b���_���a6�{��b�.��u��aB0?���\�dþ�DͺlD����/_�X��rG^f.�Bȹ����à������T ���K8�/�J���]��Z%���jjk�t��2P����J	�=�Әi:h�Z(;��i�_
����S���O��!��:��W��A=F�9J�=�_\��`�����	��l�oixpK�mi]�(�?���6�¯����	s��`�;���x\���à�b�tv��ϸ1V�r��F	n׽�sLOOܢ3:^������N�(Dܚe!\lr��H�4�3q��O&�\9��m-w��ӌ2%v�C���n=V*��� Iw�9�fj哆W���f�Bo6�]���}@e޹�4X�%�cZZZ�NK#�" ��cWRM�e���|ȑ�$e�;X���Vn>��w>�=�
B)e���pv~ q���I�q~z3��3kP����[���{�7� ]��07��AY�8y��۪\SW��kո����ANC��c��jo`P��p�'�Bo���5�/mx�_���L��w� ��ȡ��jɓ��eW�m0�&�2>wy��m��dCDj�40	"gGs1�2K��[UY;�sQ�dW&�(Q�55b��/'�������h`4�a���}� i�%��(5i'3f�z
@��_���V�(�x/ �E/����|n�7����>|;_̰6�1��]�/%����y�6X�,2�)M����|��W ��Wn�鏏�ii�|hh��ܝ�;wo[�s%�zfN�G[����~�5��Ɩ���!��K9s�\I�y��(9�H�2}]OϿN�CJ�y'���ͥI�VQ��Lr��T��Tm�����Tؒ�E=v��6n���?��O�撝v������2B���֏��������.������3ȗ��/	bΛ?���Mes\'##SO�����m;����,Qt��W�
ʝǬg�5�E���U�έb��0;!
�8@�ǍVJn�~�Wd�8·4�W��JZ!��+�am\r���xy͒Y��q,�%�U ��n�yf�Zo����sa`J��c�
o+�!�:-����I]�:��,��E/	't��d��p����g�u$Vwa/�!�Dօ:M�P]W�Q��:*���*ڄ��_��s��\t�]񇌚y���"���,r�+(o������ �x��/7�_�&q�L��acf�L�P��{󤶶6�OW���VԼ�]�t$�6����/�[޵dTW�&��WqG�j�`|ۚ�A47��ێuċ-�^�\�H��Ƣ�VS���Y�>�N�K��[���'ӃFN�$�����f�	X����o===���eb���J�_�%�
sy��G���H��1�%��.S�HT����]bTb��q�n��`C���������%J`������WWɞkn$��Q^s>���\��K����.�c��nj��k-�&K=�8�٭��@>���O۷8͏@y� G�Õ��2�ͧ�;��30��������d>�p��@�*��H�v0���	� G�lu�	+++K�
g붇��
h�z�*8K�
g���?�<'�ԿàҦ�~g+�k�!�\J�%�qb������2��˵�n(I$��3�����o��,��Gn�Ʒ�k91�MSy�A��𞔰��^I_�<ϯ��� �ÿ�f�y�[�om�@���^����}�z22KOK��� �}�s�Ƿ�r���7eetӱȕ�=\N��	_J���$:3Sf(��s9s5�K����&ݾ��z�7�W�'���-MО�<[.;w���z�wCC�; ����x��3����+��}hcQ�@����O"y������v���g@��xB�ã'-������e-- 럀�y�����t�C��6���PJ!��A ����m}		+ݸ:zu�O����� ��Ce�0Պ��8�C�̃����mzHd���
q�L�n2�x%|�	�B(_���L��BrvZ7y�tl6
��kWY+VF���YC�h����1���h�_qA�]����k���d&/f,������7��eff&��
!�v���3�V)�P�麝'��?8��0�����f؜`P|���y��ݲ��vCUm톱�r@ IC@��XM"Q�,���rx�ou�Jm��9������j�G�-���|�R.ž��6co陋�-\�z�-N�I�Ζ���bk<��&6�qu�S�0�{Hw�#$�x, )T(�/���C�\P���Z�pu��]�
SU�=[!�o������mf�sE"�H{k��ps�$0�H��p�ɼ�
BwmS5%����499I�[�k�����Ce�c���3�1N��n�+)"PЫ�[��~����Aùl(o[�gk�`�n�oU��͂2��̠j��[ ���+�����x��LЫ��jq��4�
��")N�� ��d�6�q���`1�{��y��wK�G6$ڌuO�[o�C������Ow�����z*�Z�~=v�)]���G1���Y����� 8-tn���-#3�^V!��y��C'M��y���I�b�w6�����c�/�W f^��(��]��= =�ӂ}����S��1I�g).x�u�B?זCq��N_��`q~�ܑ�u������D���������|�r��6T<r�Jo9nggg�(� }��𧷯jTt�n��T�˻�C%%�!�?-=�C"{F��&3�Z�(G�i��:�/��͏ U ҽ�����qa��������J�T�#*����+�����x5<|PMo��v�=�"�_MX�N��k�AS>kJ�¯�&Y8ly�3�E~��+�&�'�/�cZ�!�+Ռ�C xe,���

ok���iɒ!P�W��q��K�ӀB\L1�F{�`�P����)]9�'z�`�uW��M!�v}���K��<�]��~�?�2]'���z�*�_ ���Ey�°>� 9(X��k+�e!ߞ5қ��<Lq2���p�X�a:I� �gCCC@�8�������������I����*++����q�(t���j��5��\�>Q+�l�֗��b��^r�\Ay�����o�$�V"5�]WH��? 	.��
=�6�������DK������5�< eh|3º��M�e`���xc����oT�T����k}d�;<���w[��*Z� &ʷa��z$�.�� �X��M�˝K斖����H��\��0�75}��۽$��c L5�L��?y���R�Ҿm���q�����N���߭�����9e3�Z�)vh���)i�t�_Xw�&m�3��.�'��Z��N��}�ӝ�7�Q���3J�S� ���"t���R���1Ł�As��F���o^�U{�-�{�Afx`d&���,%��*�����]0�ɸ���`r���M E���J��Cr��S^�6A��Es�[{b���:�A+9ߕM�f��۫�9�X�)xLyӰl�T��h�C��s]�N\@��g���\9��tl�i��&b���ߐ吮�c�l���oq�G����|�7���OT�sMy�+��fɸ�L`�� �'�(���~�P�a�����F�&<��66Q�1�r��	��,���!��_�ٚ�J\M�y�������/Ht�&Q��<�ƈ���+'�S�H/�n(�%%s��ê?Ѕ��ޟ�Ԭ��R6X~���
I[��HY� j'�ڟ
�৫���� iu0z=�	W�!�7+�,s�����Ĝ瀽U�3�`��鱰��>����b���8���Hiz��o��Ŝ�z�))��2������ڙP�80��y��2�2�P����q�޳i_\ƿ�����mp�>|��$?����hqD����*O}��w���\�փUcB$YD�_�Ѡ����4�J5,�n���`���^�`��/��ޭlv�-R�H��ѻy��s(�l�٥z.��P���e���j2V�L���<���S�cG)NV�d9�s����-�@�;�����ݠ9�8�%�BTR�8p�D�ָ�v�L 쪔[���?�R��y��C�V�&��ըt*�s�E���_�;�+�!$��l�tκ��u�; V\ V�ίzJ�)M��1�S(O��n���T��Q��S16J)�t���ͩ0��z���~>XB��3���$G�7�[3z����`�`�<܎��!|�Z����P���������݆/ĜܺG��@zO��� O뜥L/����2aQ8�����5v�ɶǝ�nay�������	r� ���ډ�B��N��{?�I.��<o�?n	�[Мi�(vU���XC���>%�su��ᨨ��Z��,Y��M�=��J��{���t{6>yL�V�Vf�2:�ZdVXͣ��ɽ��qiL��;�����3�ie���ϩjii�[X�C�pR�Ү�@��,����w����m���,�#�� g8��s5�d��x$?Y@����:���+ɪ������ /T��ۼ�������:�R���T8�r����,)�Q�-�W�I��w�'��s��� ��s��q�#q�sQ���$�H����#����\^C����ч���(C�U�Y���m>&Q�_����A���$��~!���I���J���X��}pA-���s��)�0�
x-r�'��ά�E݆�:���Y�^���ؙ�Ѝ3؍���]����l]Z���y��27�){���Ӓѐ+i��\�����cz�b���.wy�i�SԤ}�%|����s����Z� �jD~�-W�4K���83�Bi�L��ģ�y�\�s���#��^_��#�
��HEL�"���2��DE��6[eA�'��������/h����&���A�H���S�����4{^YA~����J �`s���L��i5�I�k��r@c|D�Ow��eK}K�u���>�����E5�x�~��������^A��/���d�}HG\�p�^��=*�P%]��t����s:���&�����åi�ƚ K&P��F������&�dfʐ����wg�=��}�Y#a�]b� �acZ͢�{/hٳ��5c��gƀE�c�ɖ�A����G���^�����?���|mM�~'���^�+˩i��D�Ly_���� |�<��sM��O�[����7���N�{CM�7�b͈2�W6��$��l9dIf�T�U��2�±Bb���,d�8��q.x��z����]!�Y�?��M��Q^�}k%��er��'���L���׃+�y��G'�J;����h��b�Fn�.����*��o]@h^yV �0��=0$q�8	��^��!��K�)~��� x������N�Vv�[��[^�[��~���d�T^�l#п�,CԨ9c���%BnG�3��l<�a@�t~Ս�<z��e����郓����3�h�@��Rm�4.1]dWE���A�Q��ӒѢhÆ���W�K-��K^��(�������،u<nq��R�(-�k����wgc|I�r�ԯCF�s�lc��UL�R�mw/�~o�8h�<��'�٢ľ}g�z��m��Z�4n��<ڄ��UZZ:��*s߲���3������d�IKd�\	�[�8T��0U4�~ ߓ��[�h%����{+��^�#Vk����@rn�Y_�-r^hV�'�B��P�U�#6�D�OEz�������(�z�60��0(w97?�0���9`�MR3�>�\/:F#
�2	��ؑ(֯cddd�BQ�i�>*EL?�8T{��j��+Z��%�� �w���M����0vw�n���Oa����� �Ȯ>�2L�2�?�G����M�0�|q��g�ʲ(�Q��>J�P��Nk2;'��������)��n�nu��>���l�Ͳ�֧C$E1�ɟwW�)� �0��u��t���u�W���Geh;DsWrJg}֑Q5�㵛z�j�F��]f�F����u4dZ�)�A�K����R(���k	�H,W-oU�] �R�^�Rѽ�70�A^E���W|͓�B�U	����A﫦i�=)�b�1�0�|Q�իִ�]�N3ź	b� ��S����T����쪴	����<\�F�#�����<���(�]F
&y��2�*��OV�(Kh��X���YO´�ng�<�=�/VEդ�&W��ܼ��зo߾�u�Ea2�����/Q���^wI���~	b��`���cv�1��MSCH�"����(�z��Q�Ź�'�g�֠U'}(k���&��4��+-���8@��A������WF(��=(��|��� ~�>�H$��4��ci�%Ύ�U�t��4��*�0N���%\b �/ ��7�,h[�P��{w���K�����Y�8�Z��nk����>*�z����mT��!��aB�5 ���� j
�B���x���<� 5V")gX�$��e��=�t��f��	]�l�&D������e	������V	�]������������N�YAy�/6�W�RUJ.���c�!�j
�ͩ��wj�+���z� ��I��wf��a�{�f�KY�09�������BR����=爮K�9�$��K�5���T�&" �����:��w�J�.���7c�i���s�\�8�a�%"i����cfỐB\��w;��=��)��i%�+�:N�W��x��R��.�]e��x�%BX�t��r�k'�����sT>|�P�z-�1�D�f��~�-�����1�j��N}��P���"���G�,W�hU�e2:`\���Ŭ��֋6�+E�?JA�լ��J��	�+Č����W��sQ"Uw�B�T�.�kf�'���Ͷ�e;���_��P*t�p��D�����P"���x���3}��ok��`�U�����>$H�h���h硡��2v�0�\�(?��"���*��9L��q{BT�S�l{���47%�hg����Ы����R�t"��b
�O2C�gw%(�a�xa�%�q�iwƷ�555� �5 ��7h]���Rd��VT^z�N�~K�}�ty&C,���M���&#N��ƕ�3�n8���dQ����v��g	��Ɯ�h̙eNI��1��
�c�b����^j4�y�	��.�4�A�{[
��x����5j�����[P#�V�~�US�vFw��;������ø�Ȥ#� ����ޮ�k�~���	Y��fCn�\M$7!̟�}h�9� ��;9��].�D����5ݾ<��`dU�+ P� �T>]s��7�>���� ]G�S�h;륹>��2ԫ�̫�м������km,s�d�7�D
��=�h�Ŭ{�����ޏtCqE�S�����E����R�TO�^�'��E֨������4C#�����x�wp�X��� �2�F��q5>ܤùCѳ�neC��Cw�TË�*��H�G���hFrZ��}�0<s�����_[��Nō��7i�=���d�lz�si���9 �1Δ1K��ם,���^�a�i�.h�Ov�ҋ��+�~�-��cηЫH&���ߢq���b'1��,���}���qMMM(��O��>���&P��nL�1FQ��ɉL�*�S��*7�܎��'�{�b��P㭔� ��2�a��b<��}Ǩ��׮8�t�S�6����>�l'�o-ţBd߼979����P&��L$��kUu�4`�x�F�L��|8b�����M�ň����mld:Gw��E�y��p�O��X���G�)���>*�/Nfb�GnI����b��Ί��f�%�R:hӾ7E
�������(���`�R ����_�F-.���K7���!-ށ2�k��3�+LOȅB�����龸��F��r:|��e\K�g�>����FLT<��[�^���$DKAN��7ۨD�F3AG�;W��9B�5�<��H�.�w6=�� �[��m+��������2Eq�S���<y![��<_�p�a � �W�J�i1x0�Z��/�=��]���m�B���ظ� ґ#��:Nw*�N�sU��&d�D[H��~�eҠ�ۑ���rK����[P� 9a� &���]�G�1-�3��1l��S�>�����B�	6-����i~$��#�B�H�DAB�#<�4���s�(�	�w9�q���fq�|�i� ��j��k�����U���D�Tfa�� t�L�H���rv�y�q����\������
U)M:g�v���x]P���[��F�q�ˊU��>j�&0��^������1�6�t�~21��	4�J�Fb��%�t�ϲ�沽nU��$dI�`��#��O��������|2MMj�!�"�����վ��et��M�>��)M��Ja���Vz\��O$�}�u�L�V�-U77g��Č{�A��p���|��ݍ��b@��s�d�/��K_1˅��oSS��W�E������P,��t��+�l����g���I{n�t�S�N��&_�{�-�����c	�r��(,��rx��T�4΍�;F�z`d�� �q�����s���� l�+u��&H�v`h�e�^��t�=tV�y9�|��������
��(;�Ʀg	m�P3�y���:���'�� 맃ɐ2�1��u�F�k����W�����vc�47��2����7+���_����^z�ia��k�Z0�~k٫;%�{�:{J��i�m�/n#����%�4SN�9፦ł�{�q��s�ؚ[2:�f����G8��NO5<��;��yi����v��y������s�r@d�����Պݧ_��y�LŒq�xz��s�{Ն�q�g 2p.�Uϖ�E��f�"~���%�ی��fF
�o�$�'��E��D�U�Z����`��N�v�>�n�Q�w���o�i}3>��w�ç�3����������!�`�.0VI�!���:��Od�G
�J/�z
�פ/2��l���E�: � %%_c�o�~I���N�4D�:�����u���ZG��|(h�uTѼX0���O�ujM���j��� �={������s]D�����=�n#E����s�72Gv*�<��.Y����+��A:�\�t=�v�`��2;x�qe�BS��w=�ծ��2|y���9�}ƞ[*����cW���l��L�f;E���J6c��c�����	c$:3x��lֆz(
Y�<�����N+tWOb�����٦e�yS���%KF�k��@i��Ə�|�N0P�Ӕ&=ee��Cr>N�j�-��@���K�ɔ�W��ww6�8���(�5$���R�e�0����B^�fիz�d�d���ر\��ا;��>����:�Nms��N��̏�Sj��}Q㞓�-8�򬠉<�@U���Gd���!\%蠀�L�X8W *�߰�\�1�܇á��<v���'�	��$=���S&�"b
�X��I근[s/d��{%}LPppG��%9<��v������Mw��8�q? y����j<���������]+���߼u�1�5��ʾ�=��\w�4<�\�%O?����{�GC��c���N8��a�+若1J�R�w0���F�?�&+u/c$��1g�U�����a{�E����v�V��h�EK�C�	�nn#�y�9���r�y{uآy�KQ�[M2��~�R����ugj���+:ïX����p����Cֵ��%�[Rմ[mc#���Ȼb^r��o`��=�K�� Kx�����0L���d���R�yB����L����&���
����Y2�ea�Y轋���0&nei�j�'�M|9�kz�g���� @�a)��&���!�HA�&�,}*�t�Dy�!�-0�Dvg�ĭN亀G�nk��+�f`(���G����-��-�UϚ�.���pV��	���'�H�/]����W� I��DaM�D�h�"��6��A�#�F�b����f�f��w\S�C��M:L��(�ÃK��G�\8O��!����؍���vG�;<������jU����~�?[�������HH]�`�X2��-3eV�!B���(���k��+��ݽb��������ܒ��ϟ��D�!X�O��H2X1*Y��7��s�A����g�,��ձ����Z�@�(S�<L_#¤U����Nv�6x&���1+�c��S�^sSD��I�x����g<R�暆��?����m���k�q*/�Џ����x�5"��C*��3EL}n�uhWC/|��G�z��ꃭ71�꒳6��Q��$��y��,/�ΪhQ�ii��ZȺ��8@{�Ǝ���ǫՈ�ƾ�+�r�羗�����]�X9�G}��m�?�$�u�.[2*�j���雯��]�_��
�oyzz�x~ËM ӧ��/8h-Jo��=�l��x^���)��c����'a(p�h�χk6r��!}5�?GgneUО�"y�� ��0l������ߟ1S�̨�،=p"f���P	���ތ�4��k*̊}��� d�^�8Ē_���8io"m/ ��F���<�K^�v^����.-Ɋ���ˋ�Z�z�s�Gj2��n߽�`Y?�\�ѯ����˱����_�co/��_���gK?,���w����Y�����~7Zƪ軕K����m���U�a}�FY�M�T�Y�'op�BC���U�Q��G8)��=�i7UV �8�1['DZQ������a������~C��)�h&܋��|�)b<��T�����%�>��|(�ݯ�
�q=E�w�u��5S��%۩�#<?���R�O[ڵ)��O��|��0��z+�Z�H����ĉa��?�[������j��͒[#�gF�7En<3ҜY}NC�F�3��-��w�+�,rsH����/�o_ Y	>;:����kq:*�{*{i!P��z�0S%��t�}+�I�u�
���ݤa{bK��S槳ȇ�����Z?њ�I�d�>Q�4���z����x��b���t�2�z+��{��dr@s�ȵ���%����^0�|}<p��2L����n�#[ܭ��� ���:p��e��<=�dq�L�ã�v�I�y�?��D�|? ���x/���Qj}i9w����.K3D�1e�;���Ǽ���*+V�N�a����q\e���,7��E(�N�f��dq��D��pK�9��U(�=[���`��4�3rG�q`�U��I�
UD���8�W�L��WWV��f��j}����~U�3T�r���@ʃ��!H���g��0q)�F�Ӗ=�#�ʣ�;�|_��>�)�Z��a��>��6����m
�H��3� ��#�<�v۵�y4P��z�.o3���^�+}0���#ۖ+����v���u!�/��)*�kܔ)i�&)���:��
q��i��-����R!�>���f���Ȅ���GR�&�b� ^�)te���ł:1N¼�jx�����e�kӇ�f:�����ҧU�P��������-P�B��l�٭���+c��B`짢*��]�jy^��~i��e.e��l�r�q�òހK��&}NE;MY9 Y��"g������@���0���m�:���L�	?�WO��p�>��gj���;���m�7:x٬,i�������u��***��n�J�0m��IM��UbxECC�7+޽{7��Y���k��Uʉ-�s�5�F��R�������K������)�o�n�6�9x}���L�j�3���UbML���(#ui�_�Q5/-NE�r7P�Q&�����p�8��;s���'<8_ �9��m�>�Q�__�je����C�GjD;�56��84�y���b�D���n��pn����[�>e��a}��%H��+�s��'���/eX��=���0���9I�&iB�j[5�1��Ǜ3�(h�4r��������к�u���tH�0��ff�y��_zc��j� ��r��]��(*��xw6���w6����ī_�WI���X��kcnݽ+�������w�*�q��q�*����=����~
3�C/��)1���/
��Xݼw�,�'4X��p�9���*��������Z�$sֿ��3���/fѹ2���ԗ;^�v�dZ[�Cj��T��+|�a�(Tb��Ҭ[�_�wH^F���?W��gl���0�w N�O�������)3�ጱ������M&�9���Q�t��r#Ô����!�݅���F*���}����܃��Ŝ�)�h��gz�N��UR��_]�zڟ
�ms�9+M��1�q"V�f���D��0"1���w�'��7O|<(.�W�*X�5��m�)bE�缜�k\)���b����U���x督�m���g�P��p-���i~��f�a3%��>ha%/�y <rڶ�ۤ�#���֭B��V%|0g��!�=Szx�D,R�������,�}�s�l���TUV�X��>p�H�_'<y�d�0��&5�}�P��+�ڽ4�9@�07Y�Ԡ؟K�(��RAp��W�U��v�˝KYc�a߲�[O]�0�����	�'�o�f�Z#k��~��8&�_)�w�Fx��όU77�H3m����4�`��dh���N]YYW@��#H84
.����V%0p�Y�a�*����h6X������jy��o�eu�ʼIJ��k��`;���Jj�9��MAAA��F3��K�Ș�s��D�x���67����������2�A/�>V�����Bܻ�8�g�O�0�V9�ZU5���/��;6N�W��hD��n��b|�]�a��^�;���y�yk�A>�C�Xݪ~[%U�Q��;l��\ۈ4��=k��(m�g����[j��@�nk����$@�G�-|�����W� b��Z�#^&�3�ǹAMZ4Goseb+������� s����H����.�~�c�P��
��~畚���5M��Bl�c�ޖ���V��`K0�.`�{H����{pʹ2ɽ�r��/������8̎�Nl�m��'��E�-�yp��5g~��ę��b�������JڀM;d/-Fj�	��v�j{��p�)��9kM$�N�߬:�FrF�>{|�J�Gu:�]Z��K8�D[����U� L��˟����έ�Y�wHg|�Ocj��Ԋ$�� �
p��ƍvw����OCŏ��%�hO���Y)\��/�2�z�{��7-�<�-�Z?��a�n1��%&!l̬Vм��sI�@�����=���A�͍?^����Yn��w�Ì�܌��_W>������#�cW���wj�>�tY��R�n{�c2i���A� ����S�-��?iC~��^�P���*R��)Ҍ��G��m����30vB���ľ��RPR�Qd�UP�3���%���"��\��!�__o��@Tj�����16����H
kq�J��0������8�����q����9��^�.��BCP��F�����*�sedFAu��s���%��n��f(s	X�b^y<�:�aN��l(�s�g�h��eo!��E������vΤ��"]��p�����L��S4Կ�Җy`�wh��o:���= ��f~� ��JI�4�hLTh."p�s:p,�ri��.	d�'s��>��/\�Q��nC���Ac̙�_��}�h�M�ZF�\����0��G������[���؏ON�~>YO����Wx+�䯓i�ʭ��vj�'J�$�dd�i�v�;�{8>�5R�Y�(��b�5�5J��D�]���`Z�tt�YO7h�u���W�iCK��o%��U�a�% ��^�9��S��X����ܪ��m�Vi��(5����}!�f(�ǴѤ �D�A	���
��8wj�W���z-`_X�S�G1�����Z�F���	�S=��RH�pi�?��hPp)��ݥQ�%����O��ւ�ն�)��4��{&�B�	�F���X�M������dL�)�>1���a���w�F�-E�Ga��XdAT����A@�+lhY�$ǋ�Yi��`�nhY3�c�2����t2u�Jv�i�3@,Mm?��q���p���a��ך�� �P-W
�Y�G� ]v��`�Xu��A�&s�/w��J3�|Rŉ�y'A�TIդ`K�2v�},��Kv��{��_J+~��Ǜ�
|>)9υ����Zn���X�X�v�'���B1��"K7k{���(�m�N�����Gn������{�I#���)�ſ�f�\�7�-�f�&x<5k*s��h�%k�̣�TG�A�wZZ��������q1L
�J�ǳ�� �UR��qK۔��tR���A��Q�k��޽[�$"c䙑9=��2�~qhxQ�8@X�tT/�K"Eb�DJ5��L�κ��
<����$w=d *�o��D�*M ���j��k"� N6���V,{#�W�WW�*%~����(��}Nz��2$�#/��݊��2S2'7Yj�(�$�_�;�`��A�nSz�C]��²�`�9��k�	��X����X�{I+�-��Gn�$7�5�[<n�U���N6ec��5�[�j�6�"����b��ez8�ś�������U	����S| �azg��-	�IQ�A�������[�lz_���pA���yvr0X"�m-�vZZ6H�!���/�xY+//o��My0+���<�%�+��m?I��6����χd�ϟJO�^u(bLT{��9�04?V^��V5hǂP�پ���r%�l��2V��n�������̉�yк�8��S�)A�Y��؍�}����� \SA�<�{�"��5��Ǚ��>x�<?N���`�Sf�N�W��;^؉��e c+ӱ</M������I����Crs�W�8K�8P�����_�8�%���ޘ3�x�5Q���o��pʽ&���s�@ ��g~:-���nd�%}b0����:�G�Y2.�"�W�4���p�g@a�:<�8�OWI���;G����wB*�!�t����{f���D�ZW�wV@�QD�:-�R�Us�-��+ֵ|�����BpA�N�D]QT���J� �y�r궑M�Y�H�oE6��w�"͙i]08����ۥ�;�^@�0��?�14n4�Y p0 �@A�=(agM��������(�n
����H���3�o���i��G6�\�u���$�,�\ٛ+r��}\��!���w��*�ӭ]E~�e��R�?v���E�����b��+)"ɍ���%�>eee0�g"Nt}�V-^���e��ձ=���r�e�-�(@���g���1���_܄� �'C����^�J�5��iEin��0�l@���/�4"N�y�~$��jI�߿|��i��._��W�[�N��x�"Ź���k
}�*bz@�k����9�=�`{�^�W��x�+�f� �L9-M��N�l�j�������bk�_�ߚx��j�/�_g�S�l{��4?�u��gsn@�|6)��D�{L~���w��g� ynҦ;0R��Fn�"�E/#.��{��i$�j��x�ׁ�u��\J55��I���"/�撱5�o� �+��0g�"�����q��qU�d�@���PX?�`�My����ז�%$����%��㔵��z�4T�~��s���=9<��j���DV�Rn�sxaiIM��ح�7�@���]{8Jj��5��f�~�.-T��e/Z�xJq��Av,���ّ��Rx��X�+[��-��d�#pe�%.C��=i��z5}���f�*����#�l@*I�3y�8��tx#I˴Í|P �r�~�W
=����&�B��b�۪� ��I�T�e��>��.w~��q}��[gߪ��@���RIa�\ ��0
\���hW���ZWƵEm�|�?�&��$�!�w�pݠy��i�r��N_S=o9A�J���aw�q��]��oP��ڳ�u�Q�����D�p���^~���W
ʴ�+����A���H�1d8�yZ�`���i����#1�Jƣ���+�9(��Y���Fd��*	�N����P.;׹Fw�(�:���q �'��%X��j����1��7J0LS����DuG�YO^qG~�48�˗C��V���pf����*�(�>�>�S�.���1���*����2����0o����?ً���&�L.PU�>=P+�'�_�:�vBe-y��Q��K�m�,{H�i���{����:���M����4%v�^%�@��''I�ԷӺ�q�do�K
j�*E����Z/S:�v���_��&�����}xU&0�ГKl(}�����k����BM���`5T�`P�p,��e�8ӣL��Ź_�p���}<c�1c���<ܤ�2.z��9�]�r ���Z��jI������Ɇ}	�]Exq�>͏%�#*�[M�Z��A;��v�@�T�j���x������8�t��v&�N ��� �?p3��p&6���Sn/v(�=+������^ś
�˷�]���Q�Җ~%��n�/�s�"�;� ��c ]�=�� m!x�+�d9�����';饙=[�����٨���	�k,^I����T]�� �#�u�u�~9�%͂���f��y��hr�2�r�%��Y�*�]3ޕ	�!��O�����/lL��Z׺�!X#*3S�[�}�0��;? '���$$$�=qI_���������5�~��d��¯+�����ϐOB�Z�w1sk��9-�9X]��\��4�g<{�9�u�`�[�ꖡa�h9[ҽ���(�sP�@1�#'0W�ƚ�C��ʊ�S�G���Q@=�r�17ɂU�P�����r�Г��*�����H�0Y��s�@�������Zv�|�c��K���W����,�|��:>��KD��ש��¸/"�3A �t&�i�]nݻ��}iM4ZLQn��V�Gs�wT(����俳>[g3L�6?3Z�#67Y�ɸ7����Z�����R������.��q#�忡Yq5kia�;���0�ty$i���������|K)挴��~�H��V�H@V7}J4���L���egj@�DӰ�O�ôg�����w�����K8Ť��BH꼭
h�~>�7���_� �ި୲�qY�X�5�Z�~�t�)�5s��Q�!Hљo��(�n�#���n��=E��16�
�
��e��V[W�K+�b˟齎���yi��"�*z��+�t��J_v��~et��N@��\~O��H{�L�f�7:����ٟ%���9�ؕ���G�HLa��#���r�Tp[J�t����M:����ao_*	�]|0�tGȒV`����ˁ�5���E������Ƙ�K��3�S�n��.�W�3���g�S0��D���	澬�<V�����j2�>fN�&'��k�q�P��$�&�>��[B�tKO�}B���� �#�(v�n��^��\C�K���r},��V�P�W@��	=9�+0�	x�k	��u�o�u�c~����=m
��Z�{�U��V`g�Nw_־>��l�E��uiӬ����]Hȓ���O{o����TZ9}���Q}(-�6j��)I���dK�lF�sN�LE	u$�`D�m�))Kh�[e}�5b��~t̼���u�����沼�{��s������4mѕS"�֏o��V)���d	%VJN����b�L�����PK����m�@�S�0�mn�rJz<n��p9�ܜ�c��xP�N���{�IsFn�ǉo(�D�~�MJ�w:yo��of|0��\�J?�F��zFm���]�bC۝K���6�穞���Қz�P}c���a
�蝇�E�5�я�pְk��*w^��������D�q$�h�����Գ�7�ڀwn�����\ﳷ4�a~rP=x��v�7���
�X������Z��ћ;���!�S�r�B��n	�}P3�u�R�b��桪-u�S��s[@����^a�qګ^�����>��T$�}�#ﴥ:�Sbl��� �Ū�)��l"VF{Q>��[�c�RH��ck�O�d����Ѩz\!F���e1�[xK!SD��B<�4��K'�c*��@�>ǩ[���ř!_��x`Lz\�R;�ܠ�6�YLAm+h�Xt�¹��d��/ԝL����ce�w�0m�}�2km�<�X,�߽����D���s���#@��I�{"���篱�,�m�n���`����D�_�x����;������2T��q��`�������N��Mn�ݚ��&���6�?c:j��W�K:�h��	!���:F���"��Z�m�4����-�Xm����r�'7>͆}�G������%�.�/���;���ш�b��0�I����E
5zA;����%&n�1E"�����~��H���N�-��!��BW�����cOd���tm�.�TǙ�>}T���f�%!D4�	Z�F�4J+<��u�?ܽ��P��Tk��0@C"�5���wȢ(E��H���I��lG��_w��ٞ�yXmE�jp�нկ���98�2k���mPSz��1o�s�<z���3m!V�Fҙ�:���F���hBe��GG���ښ$��*�]DV:�fi����~aٚ��m&�魎C=����� %4��C�Kh�h�wA�iM�����7��^:�#�z�t۽����L[x�����B���H�� zF�6����I��S�� L��s�&;��\$�7��յ�3�:Zg5�K������fR���Ѥd�jh��P0`�sez�e;PIMm-�4k��<s
4g�x\�_����D�9�aDu�@	���_�ݯ��� m���g�,�2���͌���#�yI�c
��C�D/f�e�M������ ������>U�֓�9��BN����kV�W}�te��pG�p��`k.�����Ptl�t^�3?Z/�����~㴥?�C=����[���>�����n/Y�����8֥Vtoz�j�W�a�wc���-�����a�}�w#jë\$�%� g
C�mw̬����;��c�~��j���;7\�C�Î���
�t�o���|ˉ��}@�!j�FU������U�
R
>ԋu����彖?��b�^�~��I����h>��L�8=�2K�������gn�ο��ɗ��isF֋�Q�����,�(޵#�v��/��+�����$	ߴ"ô\p��G$����u�s?���V��D�-����8Q,>[~z� b��]���);J9
�8����C�{K����RS��w��;\&J �]��Z��Z���.���}u7���pI�%R�ވ��/F�2Z%F���:J{�����r��Kh��]ߐ�l�+���Q�1��yg/S��b�E�`��`��1�v	��u��I�[8
���c���ʫ�tTT/y?W����e`)C�$�J� �8�B+�	욳��� n�=�4gM����5<���B(S��x�A�w�~+F���="�g�MmB��EjOO��%m/m��2#�9�5(t*jdC��!�?��cbԉ�����lgQw�����$�g_�Ѝ>�N��L��r)�m�A��ǿ�ptq�&�G�=��L�"&L������ҁE��ab�O�H~��T@:�5A���N���B3���"Jx\����_�-���>,�����-j�BM��P����#/�|ږ�_��^N%�n���2a��5������]AJQڂt����%:�A?���Da.���'���4�P�A�x�@���{ev� �(,(l��EJo�zz��Y�N$;��/�Ŏ�5���-v���Zm �O�~e�垮��D�yy./��G�҄/�?�K+FR��]�Vo+E�t�z'X:�JB*�*�].�u6~�t;��o���h���ƪ�h�D��&��ҝ��<��"��/9��T#��� !%=}ڔbdX]~�.i��q���FQ{>zE�\K.�2���Ϩ���3�A�������2لvPF���}��#"�||"��F�X��fy�Zx��Uaݺ{� ����m7��6_Hk^���W���<͙��G�N��;�}w����B�n���ػ,+�� ��NK8^�녦����f�@�z��S��)�M�N�!=��[�)�f��'h��Yz��J�����������_G�l��� %C/ƣ�|zRRr�̈́M�(���G�㑴���굞�h�GE)��:�R[~���Pq�fvxo�'�<�
Z�t\���lP�E]��������h���/�Jpy�d�(�)#{CL��S�aZ6H��C�n��ݺ���wE��V|Y�f�D�j_qc���?�Ӂ���o�k��9
l��/(z��������V���I�^�'������GA�����L��`lP�6|?c�ʌ�hN(���5���x�~���x�2~b9T"��9=���r2a��-��'`�L|�˽���H̢�6<���o<�A* �!�ؓ�vJw�m�}���f�0C��2�̵�������V�)�71���lpPPp�yX��zq��֛���~�J���}ԝ˒��6��B��+�2(�oV��9��:��nEO�f-���H�Q+ji��8[��z�˕�4E���`��Lm��5���)�5���U� ��~ԥ��7��6�^�
B)���'t�Fw<�w�V}w]�\��xE�SP����H��p��Պ��^���������
���V����������Nta��;v}��7�w�,Z#�s��z!�#
��y�����������h����	�f�FwA�8�+Wh�Tɺ0�S����W��kh�ꝇi{xx�p��=�V�>'J�z��5�Q:r��B�|#�D�>WA��]�������}�E�h��}���0tF!zXR��;�Mr�В`���ï��@1
F�A�G.�i��	�6��J��wB%#Z�B��u.B�J��*��Ц��+�n�z��.�!�q%�R�2#Jo���c�1���D�6������8Z/�^�}8��YJ����
Rtyϫ�|�EgǢ&Yj��x30V�g:7񆊥�![��POUW]ߠ^Z����؆�~��|��޽����{E u����eՋO��e�� ���+İ����|�-u����{r�-�C�~h�1	Y#a��9�/�,���������J�`,Rs��r9ʋ��wX�ZD�9֠��N.��K4�\GG-�O��E��AfУ�w���i����/���-GN4��|�A]�h<�=��1f %��D�Z�6�EM�������݃Za�T����y�n��FG��q4��;�Ui�H��4�Q�T6�f�*y��i���B���!t�Ɗ�u��u�MˤFg���`S�`�$�(F�n�{��x��~P����QÌ���Y���V?�E���K�(�J��az���`���ς
-����(c�^=��������S�����,L�S}]j�VƓu��G�E�q��S��7�j�}�|gl�v�����d��R?�FFFZ%3u�`�mC�VA�!��Ū��c�r��e{�ꇿ�&uۗ�l���mr8fETfVD"�o��c�#���^�6�m	H�8�����jIЗ�_��Kczrg�%΢<0�<�����,�R�"���X�`y��sv�K撻u��ղD1	,�S���������+KVF�D�6ڋm�����|��z�[�]����ٲLP�Bp�镚y��b�`a�`� Y`��g��}��^&+�l����<��rN`�S_����% Tޭ3f9��p�Q#��xML�q��{�N�.���t��������!=U��S�R�׉]��Z�0�g`�@�P�=�Y��(���ɹO�nD�b�Qލ����O�}�Ơ*�U؁��qn|�(��E?AA�+f�o�:i��t���]���Tw�<�-�`tC�j����z�:���g��'�:ե��u��}U��C�Oг�~��q�&��9/r��m�����s�y�r��tK���g�S�\�����s�>�q�I����.9q��Ñ�O2m�J /����!�z͘Y�!U��o���?�Z�rCn�G��+U�.�HW��X�0 %.5��t���GNu!3�pa�ꇔ���&hjC�q���=�c��=yy���d��6�i��Sj��l����͑�ˣH=���PKxÿ3 ��e[�Λ�JV���y�ܔ	������Qr���/�J�����_�P�d*M|޷�-�Ηz���j�
��S�lQ+�O�{����Fo+����Y݂�Ktd��y'�Kd=�F'�����?��Jzg&���qpY 1K����,�����W_�zH����4�f	�5�j;I��(w���O��ξ,�uqK��Pa�S8S�U|�]rs�3�RR�T�$eq���r'�s���yv1��IImrD�C���UA-���J�ӿ ���JR4!�~#x�#�?}ٳ��=�.�|)r����Y040�<�����k���4����b�\�#�{�nHn[I|�
��y~�?;�M��M������Ӽ\7<����@��|'���z��嵮ס�j�`99��������ZR�Z�jnY��$�F���8���/�!��81Y�� �u�k���tTN=Y��x��CW����j�5�ZTqRh�eb���U�X%�J`$���=�ٟ�1��j�Վ0ܚ]�r�q���=늎���.�u^R>o�e����RqOW~#]��LyE�T���Wd��~�b�����"�za�k�����y:ق��P�tV�t���l���R��|]��>-@�T�e����&;��#�J=ÿ���j�.�q�Xz�tRW�/��	<�$�L�4�e��A�M��E�fH��e�@qL��B�v�D�@�qb�Tg9�����L��r;p��:���q%`����D�
���C��MԜ���e���*�!��/'�T����GA�Z ��ݚ�;V�׈�o����?'>��^a��E�9=~��p#Г�^��/ၾ�Q�k�~=�a�������xfhH�|N�dM��Y{~���v�����Z� {��;�R��Wݬ�z{�-o�n��O�,���"��:����lF�����FVeH$�۟Ҫ�������Q?\R/���Z�zWEV�m��~����?.�&�c�����2b���i9��=��*j	V��+���䐬n�`.N�#=��b�3MKL�H8�F����&x�JN$K	��u��LCqñkd1� _	����f�g�Q�يFvU��k��K`G�$ևݯZ;�Ր�嫗�'ܣ5꼺�~ |�����8^��$c���X���I����L'V	��v/>3�n�Ѓ�V�R��� q�
�?���8����3v��az ���I���h,�d?�'��;\�%{��iI�1��Ң �qi������8i��ո��*���x��k���Fz 9���J|�0����b�
�W����`��_�p�e�L/@^�x/VX��M�6X�p���U���(R�E^��/UK�R�� �����I{��U�PIMZ�o/^�����U[�d�Ղ��8�b���T�x�Λ1�!8���� Pp�ā?�[���W�8�X��t�8zRO���l<�I�Yv���Ƽ����H���e�t�\�D0?o͌n�(�Y�pg-f��Oك�#�O� �(U�r�����#A�rRw�eT���� <}�Z��=�@)�����9�E�S��R,K�GS���ٍg�d���ڬ�q�X���V�4�)YP����=�0|l �%�j����M|�Tv#D����hrԿ.S,�1	���6ۂW�D|b�D��߱���	a�\]�����L���>���![������x��:�e"�Ig����+V���ƴ2i�C�M.F6�`�x�wKġ�������oHrӀ��flf&�A���!R5~;�/2�6�f���Ԉ��<!��N��9�Τ�L�{��W��'paO
���;�!KL��p�!�y_�U�y��e�5m)�%gK��L��BF^�(x�x�V���_'��]Ϲ�$.��8d��4H�w��O�S6Y9e@�8+)��y��I����{�%�Z�_B��x ��07�䁇p+���4\<@O|�88߂��
7F�Ӯ�W�M+��%�H�fVΉqd�ub�!�oD6P���dur-N ti~ �X?%[\��h�d��k��H��'��g�z~�84w����Ō��8����bu�L�����d*���Ǳ(B̂��4+X2�1������|m��l1�����I-�6͋������͏Yg�,)�7�8ٖR�v��q�����ui������p�
S*.�7�F05���.��V�����5���h��]�"9�/��,��ws!Sb��g`�*TU� �	��W��Z�'�#�`��;n�^^�[����"%ٲ:�ʺ� Xd��:��x�_'vdgi	��V�	&Gi���z���W�e_�,fb-��~���2�s�T����>����K&]�b��p�i�Rl��d������'&��N��p�L]ThR��k�9�l�8����dv4>Ó,�6�6� *���f:�N$���خ[��*/bLGUǪ�DʲYӴ ���-������~�_���-�[��&|m3h@� �qQB��ę��8fɕ�0��F���@U<R���o�v9	g�5]Tf"u�����U��!8��3
��@|
J��H�$k���*��FQͯ��́��D�*�����2[o�WO"��_/sW��J�T�s��b�������&��`�e�7d��ۘmD���z"��.�=q�����o�o�k�&mN��]�jAѤe���U��;'��r>ZypD�IW%Ą��9O�T�dٟ��m	Vwٖ�dCM�I�#�C ���N-�\�/i�0[BF�+D�������El�c��� ��� *Xrִ|�.��ٽ�R��g���&�ta%��U&zUO�^e)�%��E��L/�Tw�o"���2I�\o�yCC��}���Ĺ�8q�1j����p��88Q�3L���T�p#�S`nn��l�k�˥(���l�Is���v�"7�L�F8�&��h�nn��t��j���*.�@��O��䏜m_ޮ�xx`>w�L�Q�Ŀ�IuA��VЗe&�Ga��{�-D����ݦ1�1%)0�%}LM��#���:M!��1>��զw�#ޤ�>��U��di��Ū�ݘͯ8�d�x��k��
;9Jc��� �Ω��Ji�&E�Q{�q�����%s+�o�, U^ޢ˽�}��0CtU3ׄ���I���6YM�@~y�{ǻ�Jf8�Z�\�,V��QY8)e���As�Vt���	���,�լ�����*rV入�Qug�&�������\V�e��E�brͺ�9�)�)�_����sH	Oꓹ,�0+R"K�,V���N������e�I3K�(#'���M'������Lo)�'W$�*0{V���>#lGM\Y�A{n���*���P�/��]8�ؽYm���<�Ol�utm�Q��hV �|�}��=cJzo�%uΣ�����_+����V�D�c�j��SS	�:�t`�0E���!Êam�n+��,��#K����G����FM�m�%e#qv�yq��z0�_u	!%1�"eLDA�@����O��h�8�c�J��AN�L��K>5����n�8dO H|��G���O݇�HZ��P�+@W_4f8	�����.�n-�B/���Ǳ-\4��r�S�;��\���6�-�o����ݎ��<G��.%�/?;U<�-sܴ)�Y&
���dK�*����M���Ĥ���f��� �7+�1�5ހY�l�nq4�ͭaZ�g��� �l����{��-��N�!���`e�,�<�LZ�J�zQ�o�Ƒ�~��ͼ�A��S��b������O2���`E�"}����=Ye�Gtd+?+C�T�޺�Y��EM�,SCV�u�\���,����ø���Eh���T~
�Q�٪�*a� ��tVc��2L��"=�n��0��<��F��~E��S�M\cHF�'��j�4���"f��x��d�u��u���S�H-<�ԋG�!d���#�I��+(̵;'�J*�2M�NL�c�t=�E@.A�cI�­�4o܍6�&�	��"s��9IN�m���߈�jv��FQnv��3a����df�̩�|�헷!ȡ3g�����'aZ�y8�5�`3L��y�� ��!e��;��}�+�E���1Ya��/(���\Lv6pz�]��z�G�4/�H���f�6)���Wo�,]��H�4�2�8�W�o�'�e�YU�*�u���{���ΆS�۩�ז��d�X��N4`�4�>�G�!E)D�߁�b��������Ni��x��`3�3[����|�a�.lfz0GM�o*�\Y
�	2JE�=�c�6��)OiO}=�߰��G-�#�N,���cZ�X�9?���{�'/*��_��2�L]d���B;~k�l��m!痭��CY�t_{�{�lKn`�p��Y8�����wC:Ka� ^�o�[��ךA�CHq��!�x��$��9$v���!	�����A���
�}��ig[8[�J�̏�������uQ{�ٵS��چ_?(G�����̼?C8���g]����F��ܵ@uBЧV� :lPI2;P�9���qm�:�PrVH�Zl#(�GqG5L�wJ����ag$�����,�lyr�T�3���P�.:������h��f�����/Y��2���M�}�']�d��Ւ�|�
�K��%q3��#�{����#�`�e��T�i DSM��	��d�����Þ߭?�*n�
����8d����cʙM8��1�=������2M�μ�w�_=[���9g��gc�6�Z��������E����_<�4{�-�^v�p��V9��
�%y��f��4t�~!�
��7�7c��y�\fn��Q�1�]xd��]y
�'��4�cI�mF�M+�G��fϨ��{�~�� �����[��+ᱮ��S
.Uj���H��Ҟ�`�<�j&����:���Ű��:�Шe���b�\N~n|ihX�GW���������o
��AϋƿS�p�Y�XW��Մ�]�X� z��p���,�����F#�e23<\^Z�U�P#��~f]4XgtG,�4��q�pT�TG�z�o��&0��}.�{�)�(F�b�ȓ�S��"���^�����Yb��!no��>?�7���[�!m��Y�{��BC�G�X!�Z���|��"{ZƳ�)��I��1ΏӸ�	����<�:S}T��7�%d��H���,�!b<���xϳt]��O%{��m˽�ҽ�6|b���U�o�=��v�����Vk}�]�����u���Z�G�0��H��������Yq2��vf6���Y�¤n�O�I��9&n��ٕԢZ���K��=ůw�Q� 2�O�K�︥3ИG�Y���٧���b�'h�J����6�sڵ���k���z�̜ �<������9�ZGOC��1Q�U�ʦ����n��A_?d�`�� g2G7����5���"K��ck���$p�к�G����1[vH�p2x��m�M��$�`��l<�yx���vs��5���w�_C��/����S��O�?�D��O�?�D������V��8����i��c���ʬ=�^|�·��,5a��dŞ �`�_�6����	��Ͼ���D㋶t���������m��������q���{��ה�K�PK   *��Xj���(  *  /   images/6c8b06c1-8935-4e1c-b7d7-4989f9141afd.pngm�uXTm�7:*�c�� �"C�  H�H7H��0Ð"��C��RC��tww�PC}{����s�?��{Ͻ׽z���A����<���K}x�]g��n�V^J�w�IY����z�!0���������4�@ g�ߵ)S:w��@꽨�;ts�#�Z����]'�����(1f���p�'����σ내�ߚ>��	����jy��q��l�$R�Zj]S��x��c�J��_ٚ�����ht5m��^�\:ݭ���ȳl�U98,`+v23+�ϗ��zNb?�l�#����-A��I��B�S�j׀	��;��rrr��������Y_�~�������Z��7����4-��~�9&��˽�y��9.�5SVV���k`�"��ں�dr,��VFKK�|�?�F�P�l
lm�D���l:&zwסb���ka��aa����VbRRR��IN���[t�؊ҡ����cWed�S6�-{{��8.�鞎�������VXH_b�kx�+M"�#M��?�5�C����^[M����)ZZ��G��%|QUuo�@LL��&�,�V!��Str�W���F9�:� ��:��֯�Y�^as��Ȍ�t�j=���6adZm�2���)��~c?qR��Ü�ʓ��n��9]|�/�rz���t��g������j���\:vB2`C,�����1D�N�p{d�5�C��Y/*�־�M��k>�ܢ�uW�ջr���҅�bҜ��� 5AXp����g��*�C`�x<��e�QbE{��T��`����{X�$F�
cTZ���)=��31���S��g|Kb�:PX��7L�c�t���d�#��?�@C���O-��MO�$��0�� ����	�7��m'���'LYt���F�(�,������/{g����`�m�����*�[c�%������2��b5�-J�\���z� F����>������'jĉ�#ba�|�;�=M���\9.�vt]9�k�!���Jm%�3�}����N���;�<�[ZY�������M�����Q�������uS%jy�goɣ�Ǡp����1m5T���^�ŵ��T�q96'0b*������J�SK@�u���O�~=���´��ziq)�F�Ģ���XL�,�����e������Y�^)�0���/=�=�7�+N�(~�O�L�H?{tt�ڨ�6������F���0mH�M1평mt{����Vz�������7��_r�2���!�R���"[M܏��|��lHθ'����xΔ�/��'��d�el�h�EE�靟�u�k��'^����+Oп��m����p��XX|z*� �b7Y����E�P!u�����,���Ó�,�EF��z�g�\�����n�h2�R�i���hk�b<��.��R�s��r2�x O|�؄A�E��H���<�>TEP<�Jc����������Ư�1w5`�[%?�j���ܺUc�h�����΃�:�XϜH,I�$�v�w*��`Y�tP���K��)�+* �:�H)�1���f!�J�����K�!��?����%5wT�Zrc9��)�NH�7�5ʰ4r��~F�K����X[w��J�}@JяJcI�������ʵ'^	�2T��pv��Or��ĝ��+�̜r�1�$�ldo���85t�q�Qל0��8c�99�0��#�Sŝ��{�7i�<gu��E�6��{G��!�9�/�<�C��9,,IvC�I<���ϝ��{J�g�h|R�
ޗm3I�����䟂��G ��(Lȇ�_��f�"�zz�I�.��)�O�m��-�Dt[�l�;3�F16� �g�J����nCӺvB®?���n������9
��������^t�9�9
�C��癜��5KM�򡵪ZZ�Z�;K���^�|d�_֐12
@��/�'ˣ�W���Tωh7�R�74�>��҆L_V�,��(��*���Ƕ�Y��e)���(C�O�R� ��
9Mj�X Qk09kf��Kg����u�]�QSާM�����MX�ْ5hԞ9�NpbV�wb�^��.ˎs�$���"�Z�%����}������ivZڵ#M5�[9Խ�͵���A�>�:_��q"F���{4]�[�V���?���B�;�Mu[��\�X.��r�ӗ�gY��*B�_���E���q/�����΀V�םt�I[YY�d��)K��K}k�6PD�)�qo�9o$��5�7�E|���tQ��#����(�,��c���2C�N-\3��(���{'�U���0�	�6��(.�qldۘ��>oy���4{��"����ʓ�V�d�SZSR*~)�Ɂ</-�(����ujPkؒ�8�0�4�s-W?F�w^�^'.<��U����)������[s����ʆUא��JNn�<��y�y�VH�ňU�76�G���� L���W��#u~��	�~��,������58J�搬^��Hz����<vXc�钣��Ҵ�u��ÚW�������.ѥ��UT�V#�

�~�lf�a23�����P����E�
�p�����g�g�7�k�g�1[tU�l1�_u6��ʍ�����j9Wc����\{l{��xzN�q��Vl��H�H&�>[�v�ه��;�s��1._��@[8iݰ�Eo9��5ic��#�a'm[�7�>B��^�2O��M�p�Ō�s���w�$||�cL��ΜⱿT�$�^Z�Xeܪ�y�^�!���3�axh�C�_핆k�������tl�K��]�W�>��1H.��w�4=���Q��:]���-�'�G��0W����K��]�*TH+:+s]�|GnO��f�ĝ��_�k��v��>l!�9����/��h<�&{�q�ynp�okbՍ�m���꛻)��Y8_1}�K�*��uyR?�]�[d=����Y�U�vRs�K2͜�$:`�[������1�Q��#��㲯_��F���n�������3DapQ���mcA�q�N9룿ce�oݝ3Ղ_�NM�|]�QJ�(�yq!�|W���yO�Ta=*�Y���%�4�AL"��
)~���o`���8N�����P���C��2\h�y�E߈mM�������� Nٳ���m)�`��k�ġ�!�qvڍ��܎�퐮�~�u�!�sIŢ�}(:��������<6�}�!�9�ʩ
�\1'U������E�w��p4�썖.cL ���$~��|���^���I5����.�ޏB�\�kH%�M1<bҔaf�qq����-^�z�ǀ���H�9��k-�!�]+�D�����2��y���	���a���A �Y	'�Кe���\3�� 	��!�cg�*���L�7�l,ۉț��d�Ԙ����j_�IHN���;��i�o�H��T}���z�C�NTr�T|�;�+f}9����H�3�%�.dYw�]o_�v�_$����p}�x��׍*����c�"�#G�3�x̨�5(���M�I:ò敝7���w��l��,KM��wz��s\����4�����t��]a��:�a��84va�� ;�_Hd�m �b1�Ly+{�;���|�CM;�DG��qv_�������&
��?s�I�����OR�A��ۺ���6�-8A��}�vu��@X^w�d#V 6��̣���5�	]�Aڶ'%QHYʻA�cv�u��������>�����gw�.ͨ����N���L�"-ǽ����\��)paF�0�����4 h�W�RO~Q�3i@=2�#m��?��D|��[x(-'W�W�f�'�#/-M��-\R���ϟ�2j湅C��&������,�L��f¯c�|���[wv��fb�~��J}9��[����[��y:�b_TX�r?]�7T��:�'7����!��W���z{,S�f�w����c;�~���"��6(�����[��Eٛ�}[�L�6��\e@PV���m!���^$�f��J�ۣu��zT����K_S椚�U##4�_y�̱1Z{���G��{��?z�`;���AO~�Fm�B���@?�֦�A�:�+X��k��=4�%x�~�X���Cm��޳N����y����ܼ>��1�5��e��\���@��Ġ���Թ�>�\L�*���=�0��g��@O���#"� .n�� 2�5$�{�0�B����D丁K꜡/+�����U�G%ITv�Q؃P)����x�2���yb3������{Y	��ze�߷�S֠�X�	P8g4eg�S�+V�Fa��e45�	@�^�BDj��$7(�+o�>���@$�����ZC�tmP��LQ�IA@S�e��"�x��Ҭ�E�����e�o;��h��r;���/��3��cJ""�o|j sR�Y���Y��:呅5�&���q�l��{[���b�8��m+bm�xᮡ�D����Z��Z�d��KJyE��6%@	�~z���6����T78��GPO���(��)�SU�I\\\��n�v�y�C��,� ���$�"E��uעu�,���PV��9:放�4���$����O�-ϭa*m�S>���5��W1��`'o�7�� 2�*Q��N$�&,��"I�^x�*�C���E�{Et�!}��#[��<+��h�jk�����HF�ܺ%������v+���%]dP��Y�cJ�@��W��r���,�ve��]ğө����y\@������hmm�B�v����ڡ�5�����1�њ��ĘA�B�pN��A�����)���n�>��R5��N�2qq/��"�}� �ΐ�/�o{���h17���?]w��2Y�?�Ғ���-��f��?�hO���J�/�}�a~��Ѹ �ʲ���6����}�6G[DU;���}ll^V�K�&�&�#K�v�p��=�ڄ���򂂂J�";��mDʌ�s��rg4�l��jHZ��K��0kZf�7:�{��nn�x,ҝ�_b=�)�N4%��am���(�W�}�;E���պ�o�?�ID��Oև��N���� LU��'����k��#��+e�����n�Y�؈`���d-�"��~{�{���q��Q�tÊ�l_�?��E!;�<��\Q����%B������= ~edg�!W2n�y��P<�H�sQm��:���@��-�I��YEp����mQ�ăE2��-�"Wh����:�����FB�~�� =I�{,��w˸���l?��m��:b2\3f�j�(3��(����`�/"�!PFǂZ}==3�)�H,6)2;�b�`U�͟~����+��
�=�ء��J����2���.�2( 8¼�H�������'y_�h��
j�i4Nؚ�1�T������ʍ��͊.[###yyEf��C��ʎ��gam��2�e9H���?7�vvٌ"�;K�GL�>3��w�~ռY׽�y��].�y-g�a��ʏj갱�,_��۪�=V�G�g��O+&]s���V�7�Y�M:ᓺ�{���#�2����q��u�6**օ��k��a!��?��F+��ݶ�g�M)��݈��C����#X�wzKA+��ړ�i�G��چP��!:/	�z�F4O��Z���V����Ym~a��h�v��ꆆFܷ��ɔ�ʏ1H�"���M�"��iNx�O�=ln��t��z�u<�dD��z���q�;��� I<ܽ��_OdQ�_�}��\n�+<(/7q�B�L:��al�j675��c�fqgs�-���˅"��矝��\Z �a����8�ⵗ�r�/��K�ui,���D�	TN���_t� 4.���儷zW����_Vי�+��N�\���Y|��jC���89��˞��m*�?^�*��S��$�m�	��e��q�8��l2LՂ�30�9qj���]�u�g�z���u$���ƢI3T}C	`���~�мO�-�[zz���Nȳh���u��&��D��88��"���l�I��<O����6k8�T&�2�6��Vt`h:t�w�./bj��1��(8;�ꁾ�}���Q�х�8��p]��_$�BV5����\�!!I��"N>�r�Mi�����Ŷ���~w[;:G>�Vh�����Igؾo��;כ�K��B�4��rC<�=��0\���m�_�����G����ϡv�V)L/{�k�u˅v�u^��-[��*� BB�!�����S����ݜꗯ�j��P�4�(��W^G���oj�[ם-��>��)}�H�"=��s�֭=�'B<
�bX��z<�9�q�N���#|@,D�y,���˛E�ָ���zsm.�s�M+G��J\�'��o8�=%���Z��S�=R����yb8:Io�߿�Ƕm ��_[�ow`��%���{�H>yh��;�ݚͭyX��ɪ3��k�^W�~�}��II�D:em.!O��p��>�b?NF�#>Z@��[���]i?{j��hF=���[ټu�������i�E�-�S0Q�q#3?u�q�-\���]�c��ӱ驗�Yk7��	����D�!L	�k��Jl�h���y�JIG�2����{3�KJ�Nn�X�ܳ���ly���4���	{� �%J/��?)qo��b��}�S[��ڒg�׻ ��r+����۞��'�ԋ�S͗ė��K�m���46�8�6i�٣iE.��ů��tn���yE����'��FHXC:�l��CCM�{�}OI_9���$��9!�q(w�ꊻ��{�\���-o���Q
=*��ALb�]ڊ
�/B�_TO����+��v���l���b&��w�u���Lܼ��W�Wag�q[NpN���i���V��A��X{X�r���G�s�thO�'��j?A��dJ�X�_f5l�c�Q��2zq�^'�n��66｛'#��ڶ��ν�vLl���v��{�'.)�%��߭�*����>��([�,_5�{�nD#���V%��tN�=k��ŜM[;�<qG�[�b8�-;��sD�[�b_���2�'�P٥Z����m��\�W,���{ֶz	?����,��]��_/��
��b�y���uߟL�L�K'�zGABl��ߊ~I�E���ь��S�&��W���8��*B�Ul��V���M$S ;��R)�>K����q�V�U>��ü���7o�=O��ygU�%�;|*�k_pd:�%W�@SòLFj������
Y���~��/�$a�+�}*�{6b0(t&�EL�i=�^�1.<B�����\�C�t�*�BM_e�[����@��4Avv�L�[碊���{i*Y�T�{��h~[�
�D�ݕf�������Ҩ���D�h߂��F Ovp�����sy���
�u�>�g�aa��-er"��"uj�g-��N��wɈ��޻�
���2h�e�߳v�� R���T��N(��}�ml�[z�[����y��QrE[����Ӛ��\�m��M��c��n��h�ʪX$l׾��j$;y�Z��tPI;�W.bSR&�H�����t"����S!	��mg�z�.[�1lV�%��j�{��U숎�o)V�%3L9�r�n�i�����BWT��ky;��s~�MN8�
��N"���ýϾ��y�5]��fFUlY���)Ș-[9�`(TG硧�6��J$'���Kၿ
����ذ������űu;��ݍ#��Ե:
˴������h5���K������m�XD��\/b��h�=7��c+M�r��"��NB��w`=�t^SN[���~�v�|!a}�-q�9WO!��s>��>����yH�R�Sԏ��O6�l���C�՛V)�4	ĤSz�+y �Qɛ;��h���y�y�]�}*�~���܊i��-�(̐~y�SQ�ӿ�R�x# ����i#㠞z�<��A�S�I�]Ϸ�oM�d���дtp�S��,�S�U���{Vk��r�a�>�Ps���v6��5����F����o�M���+����E����0]�)�\�lQE�ΔR5�kw�a��Ǻmk}l�|�ڭPu����d����)���V��	ŵ���w�rLt��j	/v�͖�d
�P�#�c�g�aԇ-�w�l^;�2g�W�<v��Yy�H{���JC��ɬ�Y�-�k(��)	���苊i3(� 塖���1��,�\�~�do�ۋ���� �[�&չ4H����x0��{�D"'i6�Bi��tF�5T˧n��u��{u�:롤���D�g���XV]�R��ա�r�߉���'|�ŕ^z/V�t����LMo,���v
wmau�?�8	��=r3���٧G�5��hD�샑`���f�����G9��+e-+?bV�i�@��ޮ�gDJ�I�4˲u�*��AHH�`tӹ'����yͧjX�\,�.��?J.�:�*��GFt�i�৮UKcT�.�Z��?��E.C.���v�C��
(�`cd�&_#�3�.��M�e�Y�(<\��h�Ő+}�vW��xCx;$9�S��#?�D�f��{�a�J�֓�����~�{"�G|��gZ��gPO��Sb�XZE%+IX��?8T.ۥ�VP�եo�E���ձi(��{��c!�Ƌ�T:��;;k0zL�����j�y��w�=�=���B��1�7!8���;j_9��������.��A�a��A� >�z�b�C���-׷`j,��@��<̥o���}�ϣozz��l:��5+����,��Ay�gK��=�{h���?}"c��:���k"Ŷ�w^N���vy�5W�=�k���?ٻ�^�;��)n�r�Q$ 9�H���<P�:��u/}ѵ���`ijI��g���^�ُ'���:���>Y���%�3=5��kT����������Nk3�A E�s��$ �����[�@>U�hqT"r�֢0pp)ԡ��6h������حs�`z�q�i�	 ��e���!<�>(�@o#j���*E��Q_�H��%� zP~#3-������.�(��>~c������k�������^��4"NJ�zRy��1�8Q���j�~�yu��
�(!)9	P{��Y�54��̽,=^
�sX��u�G pUUՑ^�w~���M�Y2@Ew� _ϟ��u���^�t�VH�s�s(��)����3��GWn�����Ϗ :����E�gȈ)Z�?�\В�~��b8s�!�^)�+���W�Q���95����Jzz��Gܒ�\!%�w��.�7q��1�=KKnQ�C�]{��?�� T�,�w�4{O�ɨ�IqE��9e�x���J/���I�6{�3�^�C�]�nѧ�m)m�Wj5�J�cB$�/�.�{��]W�e>��.��,,,���m��e2b�����E��ػ�*�-^}��'�%�-�qjx�2��K&��I�#ݦ�������{�t�}���å��+	W�@^��RҖ/?&�Gl
�9e֠O���Р5:$?Wr_��@ gZ��d�\�]>C��W�s���&�C������^����1r�h1�0�m0�JT
��F{���^������Z�R����i��Xs���*��*�\�h��;^3�a�%0�o)��
�<�����v�� ��9@���" ��HK��'98���(^�;���/ ss�%^"y�����y?�=���/зLFf�R��GKI0��ҝM�N~���)�?K�m�\�Β)|RH~J�J�"4TN�\��
0�
�L�U��}�;�)E��+Ek�=5�����)V%��d,�G��5�&�qCq���L��Y��f%����i��/�n��Gyf��ڜHM�Z����T���^�@���2po��J���BLAjy��h��}O�s��H�hY�8bC����`�BNZ9��#��z�@bu�{H�J�؞h�Ft5���9����M�l����>���$_�Џ6g{�s;�?NF�L$Iz�4�, p~"��F�U�R\��H�Y��p�Q������������HluE���|\:v��-\�� A�ႁG%(+)E�k�#��E-��Ec��f+@��:�P<��o��B�y����,�ʘ� ot��C��%�TA0�<M�\4��,�?�~��D���\�6��J��{Q%�cٰ��6���b��>�6����xB8�cl�W�`4>����q|��߄���u���bN��:Q-F�q�05�������
�&�EDx��q��ݡ4��Gڽr���-r�؂�����.�J�����#��o�>��Q�W	8�����{�׈JG
��>@R�������PK   ۍ�X����O  J  /   images/76768ab9-a537-485b-9af2-6ea55daf4943.pngJ��PNG

   IHDR   d   x   �W�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��	����! ��(*x߸x�ZY!Z���bY��`��TQ������h�I�w��
�( �G�QDT�A���XE6���?���y3��3��W�`�g�u��������頚���k����uuu��ZӚ5k��/��rI�d���3�:u2�����ϴjM]�tq|���s<�_|1���/��gӹs��/���?���~?��ӎ�X�u?�@f-��j�����nݺ�_�p��p| �7��K/��$�}��ש$:��/̖[n�`;�����[�|y��+W��;�5��=z�^�z��v�m��`�����O�����}��y��o��T��������_�l�o>��c?;��ׯ�����~&Tӷ�~k>��Cc����j��[o=b��6�nРAx�7�V�^�x�$)� A2�v�jv�e�����.һwos�'�C9�q��M頵�jGs|��N
��>c�g���3���?dȐ^{�U�sb- A�`��O>i���k�}��+V�0{9�쳍A���`q�.�7�h�!G�J�9�c̡�j�N�j�̙c�,Y�K��?���?��UW@`��wؐ�{ｷ�<y��޽�Y��G}d,X[���q�M�>}�J[��/k��z�-T���v��w�gϞ��s�5֎�Y�fk��Y~�k;�cq���n�zo"jj�M61�s�;Y�3ӦM3O?��Y�jU��7�܌5ʌ9���>���~��g�m����Pħ�v���b��=	1V]1�'�6���7��QY����_]�1�l�q#����2_|q���>��3s�7:�9���۽�d̞=�\w�u����QEH�\`�1w*��O6^x!|j���VJ����Q����PoG�u�������L��O3g��0Ç7�W[&����o��n�)��6�\s���K���m�ݜj�����w������b��PGMY v�o� ����=��3A7(C���!$A-J��P�����|�t�R3o�<s�G��<x�㥵Ϳ��϶?�='�3����"p<��|��`/
7շ�[�U]
<1~�&\E�*�<�t�x��n��Fm��<��	^`;_���s-Zd�<�H��pZ�^d�ö�`l+@�x���P��xI1
@аI�>)T%�H
��A�C�Zp��50H�J0���u�8ĶCl�������]XjGa�8�OT�tC8 ���w�������D ͠���S;찃9���v�m�SiYJ��s����b8�L �?��9�3L}}}_F/�N��Η������f�M7m1rQM <w�\�L� TR()�C�o`9��c�=\ �b8Ux)� �H�H�w�i'���������=�������myh@���ܨ�f�mLCC�3؅���w��}�Z�h �H��C���nu�QNjB�m9�#F�p%.�G�����A�q�	'8;D���+���BeGXZ�KeAtv�)��h��D�ƍs�GL�i�z���;�].Q������n
i�JJ
� 6;���W\�hO�����M�����#���;��SͤI�:a�p"h��CT'L�`|�A�裏:p� �E�����3r*�R$o�`��E%{��"Ƹ��;��x���o��0npp>���?�S�;@�\��<8"��6WwNv�3���p`d����Gy��$�����8q�������򜤑6�xcw���Y	���W_}�KQAE[:�F9nF�`����{衇����dD	P`�
��T��ùq��B����~,�e��:^� !	}  �^L�f��c��O�\\sK>�T�/#� ß�dD��@v���m�R���w�D5�#J�=l1yT� <4��QYM��i�mEJR�` ���B*�pCJ�
�#�TF-U4"�dh���$@ ����+1R�U����/���,���x�֧�S��V �^�"�Ρ�w��5Q|s�&�ƼV0 0 @����l��V5LjF�V�`0�� �'��q\a�sfQex��T�W��!ET&���$�!5�1�H��49��
(�¨�&I�0��J�3ޚ�'K�g�Y�9��W*�� T�T���{����$OJ�,ܧ*[��u����bʗ*A���L�<,  =B!Z�[�4�q�sc���ƶ *���* �h拳� ���l��l� �?vFu`�ͤ�#eՒ�T adQ$�K�lٲ��h~{��wwb"̦���d0�(Y�e�]AR�lJ5}jF���"��Y �(�*$��oPQ]@xX �4(&AR�n�X����AI�qfm�T[0	W�X#$�P	(�&��Zb*'Y���
 �c��bpe��R��!WD�'�R�J�s��
$\�0POT���M���8�0�~U=���j��$ 7��_�D��O�`>�]K�
yT�����ħ�m�@$Q� �����?v��kfJ����$0�L�)%0�Q��1�s��!�I�P
"�6��I�cK�A���ŵI@ 
)a�VZ�D����B�|�h3OC�eu�xVxU�AJ ��,��;b�,@� �9R��sϕ-%bQ8�<��V�w�*�ӑp�YE�H�d�Z�r�]w�< ����˾*����W�a�3~!`  K�f/e��c3h̟H��A ��6�R��L�Ȋv�ŋ7:�� BRB�3np�U(0�t��������7$b<iAE�JC������ʑid�݌$��b��2�_6ꭷɖ�������%��R� ���6%4%��^W��H�����V�kɝ�4��P��h�_Nny���5H3�ꤓNjaC����C2����s*	ɾ*n����HE��0^�O�jy��:N���-��k#�}l�hѢ�����j�H��H$�|67�7�#�Ľ�!!�L&��^Whq���Sq�4�z��1٬)�،!���%y(�"
I	�����G��PJ$R
���똮�3U`�ᗶ�L׭q� �A0�c�)	�K�x{!��#����-��PL���Gd��~�F���xSI@ ��k.�78��h7�B.� �61�CF-�W��8?�`���� �z�C� ��!��\I�ʀ8Έ'%��Jb }c���(}jC��]"�AA��_��0�q&U'Z��/IJ�Q��<G�opmar��vI��{#Q��f1Z1@4� ) "I���DI��p$*Z��9�4R�l����H~�k�TI���3���� "E�cR�:��9DJp}E�G EZ�\��Gݧ�������f�x t�v�Q$�f�B��չ�nB��|)z�
j*$;��I&��i%+�`���B"�qꀇ!.AJ(P��q�P&�X��9��g6�E��JZC�=�g�t�UV�/n�r[�$����E�����b�B.+�B"�`�rk��`>�!���!���crt�1�R.�IW�~}@��6[��L�睄\���5� 殙�`V�P졮}�4Z�GU�}r.��/q�`P}#��fz������TN�N7�vl�nݚ�xv򳒥� �Gmi/,F)���Y��/=���� �� ;)# ��l���xv�+�Dx���8a�����ڋ֧�n��QV��j���UTb0(i&<iLS`��X��4���!�B0�cr�d����lo��X�I��(�[l�5S'o�b�*J�6,_�LRWL�U»RPj㲮�	�2�T�=p�5tM��Z�^��(�=Bo*MA<)��M����a0^j
U�ݣ�
���J���>���s��!)��ğE��2�4/���+b��5�._ta�}��*WUI=P��d�H�#��
.Q�Ķ_X{�Ā���IL����_-�D$���nh�0���10�$"Řb$F}in�Dܓ�����\Ubf�����MXljfK�(�!��)x[xq*riC4���bF��h������!	�&7#/�e�>Q�=#�Paʩ �J*�l/�f��iFm�LS�?~?�
����g (LCr��l�=���Eաu\܏&�8�{Uv����(o�h��R�/�*P� 4T����Aft�Yٍ��F�5��*aRii֔�*\��DU�k}{RAs\LM��O�{�  �����0S@��&�Ǿ��Hgt
�b�*��c�'�	��ՠ�%D��T#�M�ŕA�)�Ls�)yqZs�����\�^��4Y�I0��( ����6ԗ���'i5^׬�U�Ɂǘ#)���W �R���+�����v�W􇣁���\GUukE�?y^�����ɕ�/���uӴշ*�8.�djT��N���6$�/��y|����v��4O��~٨���tJ�m<U���d�OH��P��Ƌe���f1;��50��҈f�R	�H&^!����jC� � �#�B|!��� "_�`[��Sz`䑉��/l��1>���¥��QM��D���	!��-Q��S-yC��6��@��u Rc�H�QI�h�[�t[�d�&e�Օ�x �(�A�E>���+�j���!p�iv� ԏ���`@��-m�x���_�F�eal�Z+*W�:)�>}�{%��6�{�n���72�E0W]u�yꩧZ|Gj�W��cÙg������AAKP~�嗻��c�W���I�&��� j+W���O��z뭭��	���$�/j�������+�l�Ŏ^{������M�I�k�u� ����{/j�I��Jҡ�xic!�{�Ǖ��W"_�k�(K*Dh���ex
�hR@I��� �5��C�[���kL��C�;C_YM�7��F{�T���%Tׁ���f�2�_��3S�Nu3�ѭs��� F��ݺ	�%B	�\tM;t���K�}�wRWRS��;�:��8����Q+f9:2�M#�&m�J���<��x��])��Ӈ�*`c�S�Z�<u{���RaFQ+Bs��'7�p�O�f�8@>�m���M�z�=��G��ٳ=מW�rg�8����忦����v�__���8@��dYON��M�t@�.O�����>ܴ���=�L�2%�wH�Yg���_�6L��J�jfC�Q��������m �~�]t���[�+M}cĜucc�9��t!Ӟ	�'�o���V�55f��������%� ����{?g�3r�H�����%�,���c�J0�_���@<+ڀ�M��QK,�
��*�C2f̘�oR��R�~e�6�͈���?��ZĿ���x�z|5$���O[�Dhy�@ ��{ۦ�&�T+R��m����R��~��"	;mڴ�r�z3z _r�\�R���xD��	0���Z!��� ��G�T���K���z����<��ʦ7l{<z�P��ﶍ���k;(��ӭ�� A��`ۿM�I$��}2A5Ͷ~���tP�m�'}:�{�m�l��m[�rZ��o����o�'���Of*E�ǳ	"6��j#��5�舽d&ږ#S�p�mO�v�m����؂}]�*�'O�mFOV����^('���Q�F����g�W�T���]v��&���K/��̜9�����1k��[��Ŗ���B�.�m����W�yM6�<�w��c������/���_��&?X7�w��a�W�c/��l+���B�n����ӧ� =�}��- ��!˅�r*xS�J��!���k�����M�ȏ����1�u ZcJ0h�ر�:�a:N�l��5nܸ�7�|sѩ݋��?�{��k��K�,��ځJQ&���Ǐw{BE�[f�͟?�Ύ�5l�T͛7O�[=�=�UF+�_�Y-�qo��x����A��H�Q���k���,!M�o�@�}Ujg���]�ߞ뎕KLt�W�@�a�PeP���n�f���'���?���_���<�N��wD�7���D���|F��7�2�
/FK�2�X׳Z}V��P�?GX�t��.    IEND�B`�PK   ۍ�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ۍ�X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   ۍ�X}�Ί  Q  /   images/a41c66fb-6d0b-4037-a131-23cbdfceef6f.png�WgP�i��� -�.]�@ �P���H�#�H	(B���"���	�Лt�H�T�ϛ�ss7s3��������of�&X¡���0cC�_v�_ ��8֤������)(��	J�����$0��~�((�A �"44T���;���J�I�{��6/��P��i�3}�H�(R��T��6��g�0�N���Wr�H�ZJ��HB�f!8�W8��&R�+��%�\�h�h=k�/�P�Σ�]U�����v�w�wwm�/��<�Ru�'���ik]����b%��
�\S�r n0=d;��m��S�͢ޕ	]{�2�g��%�҉��aLў$r �\�1�A��O?��vʩ{}b�~j	t�dK,�B`h-"�<��-��^�F��QUv�}lJ�,c�o7����}��r�bL����	��f���-�",��J;ㆥ%vHF��Q�E�A�ư�&��c�h�N���L�˻��~lV��f�����1Jw��K��s��jt����<�:&�2X"i*?0d���cfKZAM~��+�Jx�/˶3�Ԅژ�.�y\��h�]�i�-Otv�=W8��G��������~�&q	?=<9�C��u�a;�8�xz��Z��|�2�D?��O�)z��H�҈G��Sҝ� �G�G�f�Ϲ����`����N��9�흮�o�IlH����j�T_R �%19���TϤ��&��4�|��Dtbg(�,�WG��hu$�pI���@x��|���DA�{� ��"��2�7�r{]VX���U�^��8��U�-��#׳_�¿9(�Ef�J��M�>�0u� ��zu�Z��}Sz��{�4gm
e�f�MZyL��ف�t��Hq�z_�BD��o�F�G�4���{*|�E��-��ŗԔ70��ݢJR��s�{�2 ��#T�E~�az����k���v�K�r�y�.�0ϊ7�r�T]Y�˭�׷���8�a4��T�g]����|�y�[O	N��H���A��@�O?/+,�D���{�T"��(�a
+�w��]�F�.�x���pM6�Ͷsf�������4[��-��m���+JDƯᗬ-�7��5�g���Mtn�
���i�~�q�9�KMVZ�ϛ�����ׯ¶��2��S��j �I�וs�r�D�#Lf��������RI��r������pBE�f-��}x��@G���$���U�2Ǽ7�-�5��A��+�j�2��u,"�Z��<f&�1�
i��EU�n�ĸ�q���6�h������W�f߽�d���v����Fg��_��֢�"$���/��o��Zl��L���/��D���N�LZ�@�L}��k��>�`�u�rWU�D��r�������gHh��=��s��BJ6��)��t�k��i����RQ8d�g(d��x��3�������>?�%ᆄݦ뒖�޷��Sq]���0��샯yG��	񌵂��"&e��~��r���D��l���u��w��h�G�iR���s�y�j�w���7�ݒk�:4xC�u����TkE	{��E�smeZ���?͖��b����vu�χ�����������mMM��gyXw� �&�3G����G�8��6	��C5�<#~�&>����J��{��BD�%2�fr��6�6�T4<��2S�k�n}A���x'��r�����H�E�ݖ��շ:��]��w!��JΙ�~�.(�p�Ƈw����/�&J�By�x�̔$aeL�ܺv��խկc��L�Ć+�7��՗�X���d� ���O{���Բ���r'ٝ���#�ǯl���@b��#G��6�T�Bc��ó�C�`���7�/�+		��E?W�m �0	g�����-˲�|�/����Ã~�=�2��Ly�~��������j�Ⱦo�|�pt�ůB�a��@5TFs�����Zr#�
�����l:Q�)�/m��"��19���u�����.������������w��ʿt^~���'޸���8$��Ӛ��w��ynՅ5��Jڴ2H���Z�������6�4��W����`��I��'��[��k8%��J���q4U���G��H{�S��ԯe����8f(���7�-d�˙��d��"F�mtvx�l�@(�����RHF�@�ݶq�l>ܖ��	�It0:H��8�a4��"�Dߧ��|�o|��=9���Lc�lM� ?~���!xY$��r�¤���L~W�[W�Ė�q�y�UmU�6?�ڙM��ȫ�,h�����q�ڊ��f�A(|�����2T�F�3��7�Q�ٌR�������ᆼ����Ik���E��p	�)�����Of1,�lF�&�I�������Zz`���{qO	�3�\����^��v��{�?��k6��NK����;CZ)����Tq8@i��7*�U�gciAS����\�:��8�no����ѡtn_��Ff���ǞO�j��q��c��e���=6��!�-n�o�B��+H��u���QGEp}n��#>Z��b���z:&�H�N���Y͝�rA�H�y'�2�G;eU�N�@e��'������@�OZ�Ӎ��t�w�����v\ۧ��p���b�Ь�����詍�7�8��l���4�e)�d>�J��1��ң+�f�2\��IuLs{���ΙM�p[�ʬ����(>o��wK.�!�Ut+��!��y�3�P�H������h��ľ���������L��ͧI5/M�xW@��{q�0��:��n�o�=^�9��¬꧟)�@�)���M:;Ƽv�!���Һ �c�c�q蒓�.̣6W;]d>p�Q' @\�
�0�q�]pC�VYB�JM�28�e�6���:}�Ҵ�������~���X\�o���O�!�U�$�.-�h��7�ɪ�)-�ѯ-�[K̞�|��t�莏��ˊvQ�����r�٩�m�+�Ɠ)�'�%)\<	g��T����
��(}B�?��9m6� r�3���w�����FK;k׾��L�.ݾ��!C��ˣ���#��n���	���?mgf�0�UU"V�$JG������w�)���`�g�?�M;
��G���S���!9��g�ur�Wx���X#�ǯ�WmVoh^؂ABl�Ҭ��/��o�%h�1���0�#�*����w�X�ES��n�
�oj������5��M�/���IG���R����(3��Gd��j��^�}�V�-OOJ+!j���[��=��V}��W��4
?(�	�Pҿ����Sh���ʤ7Irz"be�m��>��=��'^m=
��i(�����X){��!�L������b��{G��� �L�:���w�����hCysX0�3���ǝ4�M^�̻���A[��#�qj#:��4[����c�vm�.a㝄�|��E�y��{&(�$x����H�ohJIM~�>��nW�����X=����������A�x������,(�r9�E�v��De��C�wE��,ŜlbT��8ϳ���5�����6Zt�"w��}1Y^;+� �4��7N�T�S/4����=��@k�,�,sgMZ<S��a �%ճh�#��̵�c2DA����N�ձ�!��ml���D�������}�
�嬠�\��>�y�B���~y<TvB� )mjB�l"��{�zL7�����f�<��}�h�&�.f����h�"|!V����	]����>8����j_��u ���Rr�M
߽>S�a�G��fG@l����nB�ʞ���H$��!�,��4��w�#�23�=@S���/?+b��%u����0�v��PK   ۍ�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ۍ�X+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK   �{�Xj���(  *  /   images/b092be47-6ed8-47c8-af5c-3a16748d9859.pngm�uXTm�7:*�c�� �"C�  H�H7H��0Ð"��C��RC��tww�PC}{����s�?��{Ͻ׽z���A����<���K}x�]g��n�V^J�w�IY����z�!0���������4�@ g�ߵ)S:w��@꽨�;ts�#�Z����]'�����(1f���p�'����σ내�ߚ>��	����jy��q��l�$R�Zj]S��x��c�J��_ٚ�����ht5m��^�\:ݭ���ȳl�U98,`+v23+�ϗ��zNb?�l�#����-A��I��B�S�j׀	��;��rrr��������Y_�~�������Z��7����4-��~�9&��˽�y��9.�5SVV���k`�"��ں�dr,��VFKK�|�?�F�P�l
lm�D���l:&zwסb���ka��aa����VbRRR��IN���[t�؊ҡ����cWed�S6�-{{��8.�鞎�������VXH_b�kx�+M"�#M��?�5�C����^[M����)ZZ��G��%|QUuo�@LL��&�,�V!��Str�W���F9�:� ��:��֯�Y�^as��Ȍ�t�j=���6adZm�2���)��~c?qR��Ü�ʓ��n��9]|�/�rz���t��g������j���\:vB2`C,�����1D�N�p{d�5�C��Y/*�־�M��k>�ܢ�uW�ջr���҅�bҜ��� 5AXp����g��*�C`�x<��e�QbE{��T��`����{X�$F�
cTZ���)=��31���S��g|Kb�:PX��7L�c�t���d�#��?�@C���O-��MO�$��0�� ����	�7��m'���'LYt���F�(�,������/{g����`�m�����*�[c�%������2��b5�-J�\���z� F����>������'jĉ�#ba�|�;�=M���\9.�vt]9�k�!���Jm%�3�}����N���;�<�[ZY�������M�����Q�������uS%jy�goɣ�Ǡp����1m5T���^�ŵ��T�q96'0b*������J�SK@�u���O�~=���´��ziq)�F�Ģ���XL�,�����e������Y�^)�0���/=�=�7�+N�(~�O�L�H?{tt�ڨ�6������F���0mH�M1평mt{����Vz�������7��_r�2���!�R���"[M܏��|��lHθ'����xΔ�/��'��d�el�h�EE�靟�u�k��'^����+Oп��m����p��XX|z*� �b7Y����E�P!u�����,���Ó�,�EF��z�g�\�����n�h2�R�i���hk�b<��.��R�s��r2�x O|�؄A�E��H���<�>TEP<�Jc����������Ư�1w5`�[%?�j���ܺUc�h�����΃�:�XϜH,I�$�v�w*��`Y�tP���K��)�+* �:�H)�1���f!�J�����K�!��?����%5wT�Zrc9��)�NH�7�5ʰ4r��~F�K����X[w��J�}@JяJcI�������ʵ'^	�2T��pv��Or��ĝ��+�̜r�1�$�ldo���85t�q�Qל0��8c�99�0��#�Sŝ��{�7i�<gu��E�6��{G��!�9�/�<�C��9,,IvC�I<���ϝ��{J�g�h|R�
ޗm3I�����䟂��G ��(Lȇ�_��f�"�zz�I�.��)�O�m��-�Dt[�l�;3�F16� �g�J����nCӺvB®?���n������9
��������^t�9�9
�C��癜��5KM�򡵪ZZ�Z�;K���^�|d�_֐12
@��/�'ˣ�W���Tωh7�R�74�>��҆L_V�,��(��*���Ƕ�Y��e)���(C�O�R� ��
9Mj�X Qk09kf��Kg����u�]�QSާM�����MX�ْ5hԞ9�NpbV�wb�^��.ˎs�$���"�Z�%����}������ivZڵ#M5�[9Խ�͵���A�>�:_��q"F���{4]�[�V���?���B�;�Mu[��\�X.��r�ӗ�gY��*B�_���E���q/�����΀V�םt�I[YY�d��)K��K}k�6PD�)�qo�9o$��5�7�E|���tQ��#����(�,��c���2C�N-\3��(���{'�U���0�	�6��(.�qldۘ��>oy���4{��"����ʓ�V�d�SZSR*~)�Ɂ</-�(����ujPkؒ�8�0�4�s-W?F�w^�^'.<��U����)������[s����ʆUא��JNn�<��y�y�VH�ňU�76�G���� L���W��#u~��	�~��,������58J�搬^��Hz����<vXc�钣��Ҵ�u��ÚW�������.ѥ��UT�V#�

�~�lf�a23�����P����E�
�p�����g�g�7�k�g�1[tU�l1�_u6��ʍ�����j9Wc����\{l{��xzN�q��Vl��H�H&�>[�v�ه��;�s��1._��@[8iݰ�Eo9��5ic��#�a'm[�7�>B��^�2O��M�p�Ō�s���w�$||�cL��ΜⱿT�$�^Z�Xeܪ�y�^�!���3�axh�C�_핆k�������tl�K��]�W�>��1H.��w�4=���Q��:]���-�'�G��0W����K��]�*TH+:+s]�|GnO��f�ĝ��_�k��v��>l!�9����/��h<�&{�q�ynp�okbՍ�m���꛻)��Y8_1}�K�*��uyR?�]�[d=����Y�U�vRs�K2͜�$:`�[������1�Q��#��㲯_��F���n�������3DapQ���mcA�q�N9룿ce�oݝ3Ղ_�NM�|]�QJ�(�yq!�|W���yO�Ta=*�Y���%�4�AL"��
)~���o`���8N�����P���C��2\h�y�E߈mM�������� Nٳ���m)�`��k�ġ�!�qvڍ��܎�퐮�~�u�!�sIŢ�}(:��������<6�}�!�9�ʩ
�\1'U������E�w��p4�썖.cL ���$~��|���^���I5����.�ޏB�\�kH%�M1<bҔaf�qq����-^�z�ǀ���H�9��k-�!�]+�D�����2��y���	���a���A �Y	'�Кe���\3�� 	��!�cg�*���L�7�l,ۉț��d�Ԙ����j_�IHN���;��i�o�H��T}���z�C�NTr�T|�;�+f}9����H�3�%�.dYw�]o_�v�_$����p}�x��׍*����c�"�#G�3�x̨�5(���M�I:ò敝7���w��l��,KM��wz��s\����4�����t��]a��:�a��84va�� ;�_Hd�m �b1�Ly+{�;���|�CM;�DG��qv_�������&
��?s�I�����OR�A��ۺ���6�-8A��}�vu��@X^w�d#V 6��̣���5�	]�Aڶ'%QHYʻA�cv�u��������>�����gw�.ͨ����N���L�"-ǽ����\��)paF�0�����4 h�W�RO~Q�3i@=2�#m��?��D|��[x(-'W�W�f�'�#/-M��-\R���ϟ�2j湅C��&������,�L��f¯c�|���[wv��fb�~��J}9��[����[��y:�b_TX�r?]�7T��:�'7����!��W���z{,S�f�w����c;�~���"��6(�����[��Eٛ�}[�L�6��\e@PV���m!���^$�f��J�ۣu��zT����K_S椚�U##4�_y�̱1Z{���G��{��?z�`;���AO~�Fm�B���@?�֦�A�:�+X��k��=4�%x�~�X���Cm��޳N����y����ܼ>��1�5��e��\���@��Ġ���Թ�>�\L�*���=�0��g��@O���#"� .n�� 2�5$�{�0�B����D丁K꜡/+�����U�G%ITv�Q؃P)����x�2���yb3������{Y	��ze�߷�S֠�X�	P8g4eg�S�+V�Fa��e45�	@�^�BDj��$7(�+o�>���@$�����ZC�tmP��LQ�IA@S�e��"�x��Ҭ�E�����e�o;��h��r;���/��3��cJ""�o|j sR�Y���Y��:呅5�&���q�l��{[���b�8��m+bm�xᮡ�D����Z��Z�d��KJyE��6%@	�~z���6����T78��GPO���(��)�SU�I\\\��n�v�y�C��,� ���$�"E��uעu�,���PV��9:放�4���$����O�-ϭa*m�S>���5��W1��`'o�7�� 2�*Q��N$�&,��"I�^x�*�C���E�{Et�!}��#[��<+��h�jk�����HF�ܺ%������v+���%]dP��Y�cJ�@��W��r���,�ve��]ğө����y\@������hmm�B�v����ڡ�5�����1�њ��ĘA�B�pN��A�����)���n�>��R5��N�2qq/��"�}� �ΐ�/�o{���h17���?]w��2Y�?�Ғ���-��f��?�hO���J�/�}�a~��Ѹ �ʲ���6����}�6G[DU;���}ll^V�K�&�&�#K�v�p��=�ڄ���򂂂J�";��mDʌ�s��rg4�l��jHZ��K��0kZf�7:�{��nn�x,ҝ�_b=�)�N4%��am���(�W�}�;E���պ�o�?�ID��Oև��N���� LU��'����k��#��+e�����n�Y�؈`���d-�"��~{�{���q��Q�tÊ�l_�?��E!;�<��\Q����%B������= ~edg�!W2n�y��P<�H�sQm��:���@��-�I��YEp����mQ�ăE2��-�"Wh����:�����FB�~�� =I�{,��w˸���l?��m��:b2\3f�j�(3��(����`�/"�!PFǂZ}==3�)�H,6)2;�b�`U�͟~����+��
�=�ء��J����2���.�2( 8¼�H�������'y_�h��
j�i4Nؚ�1�T������ʍ��͊.[###yyEf��C��ʎ��gam��2�e9H���?7�vvٌ"�;K�GL�>3��w�~ռY׽�y��].�y-g�a��ʏj갱�,_��۪�=V�G�g��O+&]s���V�7�Y�M:ᓺ�{���#�2����q��u�6**օ��k��a!��?��F+��ݶ�g�M)��݈��C����#X�wzKA+��ړ�i�G��چP��!:/	�z�F4O��Z���V����Ym~a��h�v��ꆆFܷ��ɔ�ʏ1H�"���M�"��iNx�O�=ln��t��z�u<�dD��z���q�;��� I<ܽ��_OdQ�_�}��\n�+<(/7q�B�L:��al�j675��c�fqgs�-���˅"��矝��\Z �a����8�ⵗ�r�/��K�ui,���D�	TN���_t� 4.���儷zW����_Vי�+��N�\���Y|��jC���89��˞��m*�?^�*��S��$�m�	��e��q�8��l2LՂ�30�9qj���]�u�g�z���u$���ƢI3T}C	`���~�мO�-�[zz���Nȳh���u��&��D��88��"���l�I��<O����6k8�T&�2�6��Vt`h:t�w�./bj��1��(8;�ꁾ�}���Q�х�8��p]��_$�BV5����\�!!I��"N>�r�Mi�����Ŷ���~w[;:G>�Vh�����Igؾo��;כ�K��B�4��rC<�=��0\���m�_�����G����ϡv�V)L/{�k�u˅v�u^��-[��*� BB�!�����S����ݜꗯ�j��P�4�(��W^G���oj�[ם-��>��)}�H�"=��s�֭=�'B<
�bX��z<�9�q�N���#|@,D�y,���˛E�ָ���zsm.�s�M+G��J\�'��o8�=%���Z��S�=R����yb8:Io�߿�Ƕm ��_[�ow`��%���{�H>yh��;�ݚͭyX��ɪ3��k�^W�~�}��II�D:em.!O��p��>�b?NF�#>Z@��[���]i?{j��hF=���[ټu�������i�E�-�S0Q�q#3?u�q�-\���]�c��ӱ驗�Yk7��	����D�!L	�k��Jl�h���y�JIG�2����{3�KJ�Nn�X�ܳ���ly���4���	{� �%J/��?)qo��b��}�S[��ڒg�׻ ��r+����۞��'�ԋ�S͗ė��K�m���46�8�6i�٣iE.��ů��tn���yE����'��FHXC:�l��CCM�{�}OI_9���$��9!�q(w�ꊻ��{�\���-o���Q
=*��ALb�]ڊ
�/B�_TO����+��v���l���b&��w�u���Lܼ��W�Wag�q[NpN���i���V��A��X{X�r���G�s�thO�'��j?A��dJ�X�_f5l�c�Q��2zq�^'�n��66｛'#��ڶ��ν�vLl���v��{�'.)�%��߭�*����>��([�,_5�{�nD#���V%��tN�=k��ŜM[;�<qG�[�b8�-;��sD�[�b_���2�'�P٥Z����m��\�W,���{ֶz	?����,��]��_/��
��b�y���uߟL�L�K'�zGABl��ߊ~I�E���ь��S�&��W���8��*B�Ul��V���M$S ;��R)�>K����q�V�U>��ü���7o�=O��ygU�%�;|*�k_pd:�%W�@SòLFj������
Y���~��/�$a�+�}*�{6b0(t&�EL�i=�^�1.<B�����\�C�t�*�BM_e�[����@��4Avv�L�[碊���{i*Y�T�{��h~[�
�D�ݕf�������Ҩ���D�h߂��F Ovp�����sy���
�u�>�g�aa��-er"��"uj�g-��N��wɈ��޻�
���2h�e�߳v�� R���T��N(��}�ml�[z�[����y��QrE[����Ӛ��\�m��M��c��n��h�ʪX$l׾��j$;y�Z��tPI;�W.bSR&�H�����t"����S!	��mg�z�.[�1lV�%��j�{��U숎�o)V�%3L9�r�n�i�����BWT��ky;��s~�MN8�
��N"���ýϾ��y�5]��fFUlY���)Ș-[9�`(TG硧�6��J$'���Kၿ
����ذ������űu;��ݍ#��Ե:
˴������h5���K������m�XD��\/b��h�=7��c+M�r��"��NB��w`=�t^SN[���~�v�|!a}�-q�9WO!��s>��>����yH�R�Sԏ��O6�l���C�՛V)�4	ĤSz�+y �Qɛ;��h���y�y�]�}*�~���܊i��-�(̐~y�SQ�ӿ�R�x# ����i#㠞z�<��A�S�I�]Ϸ�oM�d���дtp�S��,�S�U���{Vk��r�a�>�Ps���v6��5����F����o�M���+����E����0]�)�\�lQE�ΔR5�kw�a��Ǻmk}l�|�ڭPu����d����)���V��	ŵ���w�rLt��j	/v�͖�d
�P�#�c�g�aԇ-�w�l^;�2g�W�<v��Yy�H{���JC��ɬ�Y�-�k(��)	���苊i3(� 塖���1��,�\�~�do�ۋ���� �[�&չ4H����x0��{�D"'i6�Bi��tF�5T˧n��u��{u�:롤���D�g���XV]�R��ա�r�߉���'|�ŕ^z/V�t����LMo,���v
wmau�?�8	��=r3���٧G�5��hD�샑`���f�����G9��+e-+?bV�i�@��ޮ�gDJ�I�4˲u�*��AHH�`tӹ'����yͧjX�\,�.��?J.�:�*��GFt�i�৮UKcT�.�Z��?��E.C.���v�C��
(�`cd�&_#�3�.��M�e�Y�(<\��h�Ő+}�vW��xCx;$9�S��#?�D�f��{�a�J�֓�����~�{"�G|��gZ��gPO��Sb�XZE%+IX��?8T.ۥ�VP�եo�E���ձi(��{��c!�Ƌ�T:��;;k0zL�����j�y��w�=�=���B��1�7!8���;j_9��������.��A�a��A� >�z�b�C���-׷`j,��@��<̥o���}�ϣozz��l:��5+����,��Ay�gK��=�{h���?}"c��:���k"Ŷ�w^N���vy�5W�=�k���?ٻ�^�;��)n�r�Q$ 9�H���<P�:��u/}ѵ���`ijI��g���^�ُ'���:���>Y���%�3=5��kT����������Nk3�A E�s��$ �����[�@>U�hqT"r�֢0pp)ԡ��6h������حs�`z�q�i�	 ��e���!<�>(�@o#j���*E��Q_�H��%� zP~#3-������.�(��>~c������k�������^��4"NJ�zRy��1�8Q���j�~�yu��
�(!)9	P{��Y�54��̽,=^
�sX��u�G pUUՑ^�w~���M�Y2@Ew� _ϟ��u���^�t�VH�s�s(��)����3��GWn�����Ϗ :����E�gȈ)Z�?�\В�~��b8s�!�^)�+���W�Q���95����Jzz��Gܒ�\!%�w��.�7q��1�=KKnQ�C�]{��?�� T�,�w�4{O�ɨ�IqE��9e�x���J/���I�6{�3�^�C�]�nѧ�m)m�Wj5�J�cB$�/�.�{��]W�e>��.��,,,���m��e2b�����E��ػ�*�-^}��'�%�-�qjx�2��K&��I�#ݦ�������{�t�}���å��+	W�@^��RҖ/?&�Gl
�9e֠O���Р5:$?Wr_��@ gZ��d�\�]>C��W�s���&�C������^����1r�h1�0�m0�JT
��F{���^������Z�R����i��Xs���*��*�\�h��;^3�a�%0�o)��
�<�����v�� ��9@���" ��HK��'98���(^�;���/ ss�%^"y�����y?�=���/зLFf�R��GKI0��ҝM�N~���)�?K�m�\�Β)|RH~J�J�"4TN�\��
0�
�L�U��}�;�)E��+Ek�=5�����)V%��d,�G��5�&�qCq���L��Y��f%����i��/�n��Gyf��ڜHM�Z����T���^�@���2po��J���BLAjy��h��}O�s��H�hY�8bC����`�BNZ9��#��z�@bu�{H�J�؞h�Ft5���9����M�l����>���$_�Џ6g{�s;�?NF�L$Iz�4�, p~"��F�U�R\��H�Y��p�Q������������HluE���|\:v��-\�� A�ႁG%(+)E�k�#��E-��Ec��f+@��:�P<��o��B�y����,�ʘ� ot��C��%�TA0�<M�\4��,�?�~��D���\�6��J��{Q%�cٰ��6���b��>�6����xB8�cl�W�`4>����q|��߄���u���bN��:Q-F�q�05�������
�&�EDx��q��ݡ4��Gڽr���-r�؂�����.�J�����#��o�>��Q�W	8�����{�׈JG
��>@R�������PK   ۍ�XᎩ���  � /   images/b3182cb6-763b-4979-9bf3-a9ce9c9d7585.png�i4�]�7�V{�j���*�Rs�*JIt�jnJm�\�,bh)U��Y��J�$T����PB�SHbJ������������z����keeX�{��g�g�}�ɻ������  �� �' ���Y�b�byf���v�뾖1C�X^F1��qd�  ��N|s46b�x�[㩷�����sO[����������sw[7O�L�* p��~��?km�񒖾H[�������}�*ߤT�S����/[=eu���E�B^���G��;ֿ�C].��9�����z�b���s���M�:�B�hHr�����O�Z�V�z|���⮭��w^�/y�8��v� �������-�L�_�'�K(s��ۙ�����>��Eg�+�^�|�;�P Ik�4� ,������9�z�ú���ב[�MJ��κ�SՆjL`bP!��/���R������C��!GCU��L�J q\�د�Q���БsM��R'���P���5NN���G�D@�p7z-���l�QZue]�a���n�1h'N�<d��om��)�^�$m�p"y���gW�2{h�25�&L���ֿ?}U���~�nG���6��tI�8W���DO�V$S[�jQ�=�#��*!Y&K��B!qO��-:�|���^hI T�Ֆ��k��N�7g��6�R���n�VUv�G7�Hpy�h7Iv\��N�N�<=^~��b��T�jq�%5�&%�H��R)��(�6�9���:6�@��	�mI�������y�.?��Ӆ0 ��c�����O��;阱�%I�F/�h���ͨe-�A�5��Ĺ@�Ft5�+��-�h�R��,胏��|k�:�Vd�ǝ-���w� 	�s{m^3
��b|�ln���ж�~��o'��6�����WQk���o��҄
�&Q:J�R<HcA*�A�9b���,��xb�1Ж�w�6� �̾I~�[�"��1P��_�ugS}@�$��]ݩ����K��Z�N�1t��e��|��?��Q�΃3
f���&�P�6VH�F�7�w1/f���~ξ���m��;;�HI/k�n��{�J�H��.K�N\~��W�_��#C�j̱M�����*�z����InRU+�^5_iZ�7�0]i����5�^"�z��=T��H�T��x�����?�z@�+,�[9	�5�h�t&���=|h�8T�pz=5q���yui��
�NhL�l�0]t����
���4k�0?V�_T���O �͆M0����q{�7JO��K�%o	��n�>*9D������� Y�H�L��C���Ԛ�����ڧ�~ӑ�+ʰCm����EgO$d�k����s)�_�/h�XBٶ��i�0 �����[��qŔ8�����N�\p��[>�h�`�ާ��Z[��_��5�r*��r�执�2�����Rs��[G(�@�����@���f�&�MB�c&?�
�w�{���q1����hWs�3TO�]���4��G4Hw����ZR ~����a&���̤( �_�_�v<�Y�Q+�~f���',����[��Q1K.����ʾםI_���ב.В�뚁�'���[Akj�I�{	Y�_u�5e�Y#8��Xƪ�A�7ڽ��7i]ocA��@ۭ5d+l��p��mn�|�J�e���%��o������;����!���5��=� q�Lã�0N���d��N�sn/�2��Q$�J�aG����$��cÕ�:o@\Y8���FN��:9Q<�}ζ�Me5���x�|����E=���)�dd��a,2����SW�p�l&�uhl,�*l֚�:j�bSNygRv4�PS^:�v�ڬ �����'�Äkǻ7�I��MR���N���,)Iva{µSw'���.�j4.K����-�t/2��u�[�CL2�x��ڭg��X��^fV_[��F̈�3���N�����YntѦ�4&��$��Ze.R�U��7�7I���BG1OY�!aa��ݏUuk]��H�~@6�M&�ԧ�D諹��7��WX .�/�{�������O v����N Q�;�S`� /�Z���y�5���Hҗ-_35)����NLYZ��H24z��i��%�_�"Zu�h+��� �|�N����>R�)������ݵ��"+�4p<���r}!2<bQ�P�t�p[ev��u0�u����u�
�<�%k����~�|)�vp��8X��):ȱ�ʼ ��+M(��弨:���dNՔ��s �8`|8F/GX�/gz>"���7�B�a�/�[��j�e�:[��o��9�����<�V��}i������ݯ=���D�f��rSi��o%����ф�3�P?�پd�l����9;���4?�%��`�6>�~=�c���`�� :u,�6{�p��]�N���M3�5�1X�o�th�R+P��R��v���g�a�M[�䁡�(���g�Α$0�(#ٶ�=79��(P>	Ysf���o���J�Bͻ4��B���9�;�@�y�y�a5�r]�-ul��5���The���v��ۉ'�6�G�	q��ϧb>����L�����K�u�;�1xva* �Z-�L	�L.��v����:w� h�;V��ꇟ�>o� �[v���EW�m[�6K���k�_�v=#�������T'/Q�)&�,�4ۻ��M��H�,��J�X1�<�V>0�N�<,��@���^ݩx��f�іȏ�p��:y��*0�lqJ?knY|дn�Y��Ja ֓���,5\Q�c{���2D�4R�~�|�eM�?�«ڎ+kL�iBg��h�n.ik9Q�7��2"���%�`�*�bjN΋<��4$?!;ds&^f����j
�����r�MZ�:#A�
3p�F&��n�X�7|zw�
W t���+Ȳ�A���
�&JW��ʄ ���B��f*�,7��*i:�Zn��d�N��!�j��r�E�3`LD阜��ӽ�ӂ�����L��Т�	�T츕���U��n��sF�;#GJ���RR5s
h��YGC=�=����ܜ�<�>\�	f-�0���۷ZY�������=Z�cxp+�ܠXG8}�����^�%�I�Zd����K��0p7�N
)�XD���Հ �K�|ׯ��Yқ�V��Ͻ�v�"���&�>u�Ny��S�d�_f�����g����qtU�l�hM�W,�=f,�L�i˞z�R��>��4����H�ilƉ�� {�5�W.��=
~�>����uR_q�����kH-�K��[���ۜ$��ck4�6�e�	>��<Z�d�\'�Z|�E�O.������;V6�Ȩ� ����Q�B)���MH=�E�٩V^�� ���3����S�j(���/��ѐ��J�@�ȑE7�'����6Կ�<�ɾr(�3�Z�/����l[
6��(�W����ĉusO[���_�N��������H=9���P{F=�U0PR�[�r�jh�� ��������2ٌ=�q�?�G�[K��ţ0y�Gf��hȮ2��-5�v�WG֠"f7�v��mF_� �d�qU�VN�*��ed:�t�����ښ�t���Ԍ��s累PX#��d,���t� <`��Q����D�IˍβR�yԅ���1�5ww�9�������gI���Z�����\���ΨХc��>�K�},f�n��9ZÅM�:��v�2܎�ao���(�^��u�v����Ft�+�8䀷��������vF]0X��N���Hrf�(2A�|`�|�W¥�5)�ܺ�9:���� �;�3�N�mFb�0i*)H#X�Q�b���Sy��>5�r��n&d䓵~�ۣW�.��K>�}�_5�n��}Q}�2��BӜ��5p�`�ԇ�a�m��n�jR]��^�|��������A��C�K!y����+�G�Bi��awf���4	f=�S��Z��g���6:�s����6]vs��P�v3#����>:�15��^	�T�Z�jQw6r�8!/�a�ob8�A�pv�jtfF��(}�5��#�ku�3��)9����@~�� *W��B0X��"�1�T��6E^m wT��P�����V�6�Y�:�M��~l�D���*�+r�z����=�o��b`��u6%��*1[i{T.y����@]����c�y۔�O�M��q}"@�4�}�=n�օi��t=-��b��-��ɑ� s�����E���9z���U�։����D��$Jm��=B�L���rKq�2[�c�����C�tFt/���1������������mԴ��K�����)66�#�g���yBy\��	r\R�4��W�2.?�3��걹��e�
w��Ar�	"�m�B��}��VuH����j������]����NN{�b�6*�&Doz�ޒ��o�B��޵�3Ϥ�"��q�����TD�	��\Hn.Eӌ#%O?�w�)Y2�kX2��=�9K#MB��K��@)Ҟ m�^�o�k���@ы�W�T���gÄ�+,JL��C�x?ydЇjA͢�?7{|�n�g��i6>�7=�@��H����-����n�mB��oRR�n�(?���!>��'��0�ug�`}2{��l2&����c#����z�c�U�)��w�4���tU�E��L����R�Ir�%����r�"6q�Z>���<��ݬU���)^�3Rw�bP"���G�%�|��mX�)��Z2D��6�C溴�V�#�R6B�$¶�q�i���4ބ�Z���T�R�e�[rb���=[�b��D��W1�Uӑ�	I� V���CkO��7���Ĺ�ޘĎ�́�Y�AZ���U�8���j���_� ����Ii���1�g��N;N]�C�d��#��ŋ>��/j�d�9O�#�Hz����������?�z������My��ﺢvo��g���>�A�$�ݚ9��[�o���~��7b���F��F�U���}^�]�t@ii޾�	)�K9��r�R5�w�~�"��"4����[3�)v�
�$VK��*I��y�|�S��~��N�-� :{���eT_�Z��t�`aT��|�no�=˴�=F�n}��<�LuCp����S1�zfn?����1I���˹%�,������ہ����t�8=<��gcn)}ڭ>B��eDR*Nn�8м�[/M���qk�^0댰�������)]�}M׶��w��9���GE�E��FȣO�@�G�d�OhnӒ�eS�)����w�q.I����6�ۋ>n��;����ǳ�5Ul����p	q��'�-!8W�om�:m�w��ʩ'B��Ue.b������\��:�ѹo�Q��FӼ�������uJ�"��{<�A��o�"G.%"nv��k�Z�Z�Z]��7_*B��bc�*KG����js����@����T��T}���5��ͩx<-mfQ�MW^p�)Y��k��Ȟ=k���T���H��q���zLJB1w��'쥖~�'��^~��&߽��Mm�,\���H5��SZ���j��Y[i^�"�z��ıcB`hܾ|��E���>ά!k�%�Zsz�K�9-_c���m��?���L�	����*�SOv��;譂�\?��_7S�/��\�'�Y��JU>��ok�Du��(�f��U1�3��I�|_wE��T����@��k�yF���U���h��eo�*�* IA3�3�x�K'�o�1��[3��RV>A�M�gož	���&�-��T�#p�i�P��H�K;��:��u����fB{�m�y�����ݖ}�� \z�E�r��������(��w���V mGs��}�������;j=�W�ʈ9:���`a��<�������w7�N@�4]�޿�H�9���lbg0#*0$,ӣ5��]��}�D|�C@˩�>��O��	�D`���vD	 �Fq4&�qu7�qC>q
a�$���J��ۑ����T�I��r�}�X�'�lP�ww���Z�:�8mM��ȆHL/I�5p�}P|8�<���cm|M<�U]��o$�@���52[\��97�1��<��)���-����f6���_�_�r���*==�x����}�H*Xs�6�.'~�|�PBX+}�ۦ1��-7����|販�x� iL�Ut�y�I��ԭ=hm2Ax�+���[�8��� ���.�v�e��"�^�BgtO-�,��5���|b,\R�d�S�����;{@tU@� ET�tQ�+5
�-U�SY��c���})�j�=e��Yo��h���WȺ���٤��߹��ZO%�f�B�癲��^,yc>�2�\A�D��M�ٵ�քт}�3�y2%/����qZwV�&=Z�����%�>�M�MJ�Z�J>�u._V��T������Py���sm��NYt���t�T}dS�.$��܌&;R�\�i�d���9��7n<>8�ŷ�_��� 	~.���x[�wKb��
Fdf|j�X�dZo��d�|:=]�H���C�&��K��XR�Z� �~gQ^/��4��˹ʠ����{I4Å�/E�g��)���I�((��@��ba�T�m-�DsϜn+�[�B�Ы�\|���\_�ڞ��$�/lY��Ȣ�b�������E�q���\s'�zsIĽ��K����u�g�;��4Ӆ��n��f�	��f�N]a~?�@�zIw�nM���p#���z��-��m���9`ļ:F�]�=��KE��Lc�ޠ�>u�0�'�Բ	w0�͘�Gg��ܯ;U�u�n��Ҭs]�a���Ǐp/I�w�<H�P���V���&4�ҽ�������9O;HZ�!c��c�	�����W(h�o��̗�*��>�]�"s�lM�f�:�+��
�	��**x�_��ב�96�Ҡ��f���D�<��!z�Ŕd<� ӗ�{�ϳX\8Ej�5���vH�h9jJ
I�ڧ^���~ޞ�0��Z���c��.���<�fD��b��P����o��U���)�ͤ�, �.��|���>�p���wM���Dr��:&�b��H^A��B�F��b��Hh�`��x�yb�B�@�#_+C��}����ɤޭxК���3CI�T.�EGY)��v��0��������`�~�|µ�>��ț1�!W��L+ڦ���㇂�&|�8Xe�;̍�2T�`��BA��rA�A��|��/���ˆ��*t0Z7"{�%k�\n�Zxn�l�+	����ts��>A&��1~�յ��R��,:���;������	 �_�|.�$0��c��B�m*7�hl>Y��`@r;�x��o�|@&��웪�	)_���闞S�Ū�#�>\�w1���ыݾ�7�	�!.Mvj2Mk֩��|3I��Gw6�yS*���l>y(����/c'	��?�6E��?�AAU�����/�m΢klRJ�3�J$��A� �7�Bmc"t5�`n�ntw��b�����(<\8L?���}2I�d�(SXw�6q�@�u�.m�,��2���V�+��ԕ7V�;�:rt]K�Kr��m%^�5�|�6�幈���Q�p����.�W5�Ln�hך5e�T98N!˓ �MK����d����N<:�#�8*���0,N��F�'�f9@pG������A����1ɜ;��K&*d����h�_q�z�*�]�U�m=(�U�dx��E���Hx����D�Kv���{�Q��M��[/L7��:��j���`�Jh5j�dH MM����Ŵ��J�����;%�����4�Jؙ�A�$� i�6&�%q���{��ՙ<�͗,[�J9m@�C�X�����#��	Y��~��=��8b-�e��{��½��A6Hޏ�:<o���Ɏ���ݓl��mR���_�zn��f>N5�q�'��u)�(x��O0	��h�Ǌ��޺ᖸyP�Ҝr@AѳOi@�`Ae��������-��5��ߋ�68��O�K�>���h��)J����P��6X��}�q?���'��m�o��e�]0�>�m�*so�e7H��9�Ҁ�B8R��6�n�}�c@l%nn�J�i�^f���j]=�U"�a�R#�P�b��6j]s}Pz�=�R��Q�'ƍ��Ú�@�ު���\8۳����w����/���d�X�L�CMu�+���,�T��Rz?�8��<�����6���;�L�������"���[��u:�,����q�����^ԣҁ��q֢ �q+z�+M���|�9�[ςE�������.[��g�[�NM�G��o��%BX��	�D�t��l�r�~KӦ��W	���k�k?�̏�H����*�<�]-݆Ub�>(7A3/��cZ^�|,�>��o���nj+�!Yx�t��V�O+P��(�������r�g�\�Qqjn��w� ��,7Rx���l�yr8"�X�עY,��"o3���Z���G�3Rj��m�s�k~;�Ӥ��~}�q����f������gj*��V�k|��)��]ѵ:��N�����DGa�1�X&Zy�k��X��i4p_V�H*ͨ����Z�h˦^�戼X����Ai�Cdh�6ÌP�+v�~&��a*�����%�:�����/��2B?�ͥ�5�:�[h-�)Q�R��.���)7�VO}2�Y�K\�N�:;q�+�[��5�9�rx�u�U^q_�=p[	n�u��ٝ�)O9�'=�i�;�(1��k�֔\Dt��Wx�/\<���?:�"�<��oMJ;�b���0�DR^�C�ߝ��C�/�m�0H�K��c_���#��+�<�B�W���O圗�,_؊IR�J�~u�
/6Zs�	�2�i�(/�Ւ.��QRQ�n�I�E�ν�j���Z���t�'�]n+/��p�_�,,y�]�O�
�J����N��O@MZU���t"��t����5�7�v�w�
`�@�f+Bn(�R�R�����/ýpiNS�c�e�5����!BPޫ�ֳ�V�%�����;x�������-���[�4���5��:ёo=s���u�j�UE�k3�HOZ|F�ξ��	��I��s8�.Ԛ(��D:V=!��RD? � �깹m6q��{r��3�/���J��E��Y��Fĝ�Y��WN8��^�^��C�S����YUmv�f{9�+qr6Z���g�N�5�E���R�:���xx���x{����눷�����_b���_��&��f� �5Z1?I����a�sq�<W�X��w�B9U��	4���/��0k.�i�_��$�#h�j���{Q>�=c�	+y7v�'�������W��Y;��g��2�kQ�[7>$_PEЉĻA�ZK=����X�^7��'Μ�G��MSeh9�Q��N�f�@��dT�VkR�x�}m��q��:��l����2j���X��2w�4w�,|%Oob�>���IȂg���O��X�{�W�^R#pk�ƾ�/�y?�,�rX3�@�O�r����ք�%;Ygf8*	�>�n� �/K�%��j��~�s���Ŀ��ݓ�~z0�f��p?�'}��9�8(��`!����n��z�*%¤���s؎�C���͟�'%ؖ?�t��4�ŅUO����?A˥&�
��c�����}��ōth�-���P�S�4ZE�~��,�P��٘�u;�,U�R����y���d�O���w����##���J!~��a��	�O�S�i*�5pUxh�K�R��3����(�0�}�Or�KkJ}��׈|s�G̤�9O� �΂�JF�ŝ�T0�p��^W=��|�tlT_�7�d�����������ȿa�+���j�q�m��Yw���'l���ro��<�B��x� ��҉"��<D�P�d�Q*F�����@X���x�	b��SrRFW��5�5ELk�n��i?>���Y@7*}��f�㧦m{�5�x$�I��kz�.~������ۺ���Ӓ���<@����S����js߰*�]n'bXϓ�62�-��o��z-�oK��'p40�~��2{s&'a����Z�H��έ���AI��7�e�ڟ;#�x���������O/Br��_��<�$`�9TI�k�c	N�zxMr�#\�K��}͇;y�	N����3�5����f`���w�Ws��K$EȹN�\s9�H��mJ�6D��>\�M���$�]#��l}�L�O���p�e�&w�O��l���m���fw�/���O�"� ߿�Tn���(�;�5���������~ �C˕�B��h�o~�K31d�%����79#���"(!q���I�	��~#�*I��X:I]�R� )�����q�5'�_�g|Ό�/�O��G��C�}���RJ�m��a��Ao~���x�qw�Z���OI��)��t+����
��/�s����əgl[�.��&m�O�m��X��5�r|:4��߂d�a9�7�Z�w�����S�@�)��c��$�g��V��n�$	e9zR�xxc�r�,���5@�:�#L�?2�YNcI�M��Q,�F2�F��_ �����b2���.�/���k����[�j�(�{��MN��v�J�K&_�ёk(=����_?�4���$�r��ޭ~MI���^����[X��^�;}@�:s<���a��.�):��v*�(��:�B�0S� �^����Ǹ̵��t�����^`�'H���"�<n p�}7��a\Pl��'��O:�WK�6GC
b~�-;)���)����6�Ѱ��Fb�-��x+��ĚW�	U�S{k/�G�q컭 'R���echd#�lt@����K�a@�}�\g��&��&��W<ћ+������;�3�.Æ"��B��w��x)G�a����-⌟[���1��آ�������g}x1�a�.ҝ]9O:#��P�~�AP��􂀕 ����VF���"ƕI�_�[��iy]��8J(����V�	^5��"S��L,N9r�ʜ��P��"V�%w �upOrz�pͥĢ�A�}K��1T��!�E7����ʑhώ�=��s���2�Ā$��c�����,3��0�_&����r�F�����J����g�P3yn�}K?rG��β��+ �/NdKD�#'W�q-b�ܘ�&������� ��;2�V�S
��+��$�jF�8o�R^���v�\�+'y e98^`%[	��E=�R�0���d�Q'm)6�Z�Y_^���q���X�mk��<N���Bc{����t�`�5ț��5�5?]��)6��z�/In�_~�Tw�cy�/vi�|��k�ק�c�����6r|���*_c7]�G�]9=��0�L��%W�Z�X7�L@�+ew}�����mp���L�$�<�s\��8�7jr�|C��ݟu`���5��`+c�Q{p<������NiJ�*h�������HY�2��d}����ɦ%|��:H�"���Q�Ь�A6Y�夕�3]$�k�@��68
�k�s�.��)����R'�<TaI��*ւъ�uU����`v��w�Ip��i�s��!��z�	����%m*M�������pHww�m�a��)B�Ia�N�ڽ��KȌ�H�xZQ4/��S*Ӻ}�c��?�j��§&��t�`��A�p���1��4��"a$͚�����q�-���8���˒���9�oi���a�>!"{�q6��E����t�m�M &�&\UV�6����1���?o|t��zhoSq���q�m���ڔ���~�8+�=a������J��ΛHay��ˉk$�^����8��HS���n�u�c�4���>�^��|r~� �g%rMو4���:���"��J�Q�Zx�lj+(��:}����@�o��?v����iq�����%F%(��p�����P0m+:����f�(��J��QH�Y����U�K�1�rB)���~?b��(s�����N�ȱq�t�ⶈ
�s����B��UV�n�%�sE�!�����Y� +�0�`�w�����Ӣ)r�{nyT_�SB�'�J��-(JW�H��Ԭ�66acf8�J�'����K
R q�{ެ�8�bkt�S1�i*6����]�:�+ˀ&�1�J^�Ӝ&�̓�v�ct�RS���jeY���Vf����/����gၭG�]�At����ctz�(vD�i�c���-U$����M�y��3����"Z�_��ϭ����8m�Ҝ3(_#��7[���+��5�'G�~}��&H�t)��(�Х:���Eo����1;Ux�fyUO;��Q��VR�Ȱ��_X�e�{%f���F�T�ٍ��N�2㪥U�ʽ�i���3�LI�L]3��dŝ��竽ٳݘ�HYP����'���к���3K �b�?S��-��+��,�=��+,���H��w�n��'�5#�ݙߚ\��x՗�R� ��o�?DǤhm��:$�D(ޚ(}�G4D�"
�:�%˒�2��`M��?�T�;�6A!�����k%��kK�e�� d(�hm�%H��H�mB8nF3R\W�㶞۞�+\�A;-`��5u}��)E�I���`z���ī�I��>�*C�T k���!d{DQN����/�A�7�����]�/&?��'���vk��j&=���GU&,'��Γv��.��}z�h&�P�#���_r>�~Ae�`:'�}�#r�D�0��J��ĸ�8���^%RƤ����LH���Q��0�fEbf��#kXf�R��u�[�h���uK���i_egX�K#)N�{�:6�/��r	Bn@@k��`���.��}� "^�5k˓� Jt�����cz���9W��7x�olw_�24�>�uQm�u'��^]s���@��mWb�/X�蹃�'�f�"��{Y_�)�~��6�"�w���1�\�vCt��?�7�p=�d30�G�^���Z�Y�z ���Òy�04/�v������M�f8p�vEϚGO@P�#���/� m:��A3���_�&����C{^��$��p����,g���m�O�#b���1�ջLgp��V�"���ҫ1_+� �kΏV|��P�j���Ȇ���Jܚ%Yz������^��$�ޘ���ښ W�k���p���9m'{����6���k��Z���e�اdФF6���)f�o�,7����)��!%闌��{?��T��i����a�[.�
=�`�^���6*�&�r��6�h��>����|��_���B���2�uo�� X]�u���{{�<[@ʇ�:�	M$��Ul�T����sWë�{��OI�Hה�N�E�����w���3U��RHY*2q������@�ҋn�[��2r��zm8]�F�ꛦ�,˻d��|���3<ô�FJ��8Eè��1d�ɭV�`+��H.���nEۛ�v#J�sO�/���#@�R���@^�&%�^��iP+�}��F�M�����/8TV"mGx�>n�X�<)e_M��	�����7ˀ��;���J�x�dh?!*��"�N�Y�+5"X�xutF�@�C��G,�^�%ԪG�Ϸ��Y� �堩�,���=E�S	��}�+�!�������vJ#
9��V����/Y.�����'P](ZG#�$��K���ȅ!�0D�����-K��
���m{B��ēO�	z=�%R�jGW/���gZ�e#b���Y�O�O���ċQ�O�<��N��Y���9���n+���ֽ��$�K+�ߓ�����l-"��^}4����[����MM��,¥ؒ"| ۤ�q��O��a*�'�;�a*O����rNd?b��x����������O~㕿P����ݠ`i|i�R�o��B�����R���c����P^��l���?[1�0�_蒹���WM|��o��O?@w��VP[�t�p �p�_�K�$�y��A�����$����x3��y�w�ˀE�,NI��΢u�;�S\�G�Ŭ�H���@j�%Tݹ?C�bȧ��8U�`[[��O��os]u��_E7�ֈ���f����'���%K*�'���
�/��,qd���\(ɯ.U���Q�|6_%��i�P�.A�,,� ����ѝ�ނ�YwA�U�x8�9)#�����{W�����ھ�?�l�3��sE���x9��.ch|�?�G(N�%s�����j��M��7*�dp�&��~e�΃^��v!���~�?�rl\ܽ�aֳi��W$�+B��&1�o�|!���O��颢�|L��1�>ѐ���"��ȳ3�U/DS
�~Aܰ.u�Y�"����ɷS|o|�}������}s������+�+�ok�L��������_�r�l>	��(ҾTy3�����پw��\Tv*���N4�Wt��'� �[����'�.cx�ZO�l���h����*����`� ��,��6_-�;z#}J���|f����\�9�|��&@����6"�\���8��9���y ����F��?LnMm?��͝ݏ=��T?R8=�a�6���]���)��Z}��]e��G�5-H���ʫ-e���4a�0<�P~������0H�u��]�B�5�������	�|�s��r\�? {��g����ҤY왅w6C�n�z�9�5wM�u��IJ>���2}4�X!�D��%0Mi�u�˃r��z�04�V�m�|���$
��#�r��rQ�'��ܺ�w�;�4�Im����+'�qs�^��j^+���i�����q}KPp��W�}P�B�+���:W`�(J(��,�g��{��j�~��w�{\s�|���"��d�2\	���l�.���c��D�jҔJ�q�R]?���b�ۺ9.�hd1knY�����Q�K�r�����[�z�w�᎒%��	Ē�G����Lp�T�V��Y��Е;z����;pG�A|�bN��l�y��b�,겻��?��/n�R�?��Q�+,��ʿ��	&?���OW��I�S�&���ѷ�a*�yr��w��<�w�/�������s�������J�����ҏ��O�m��X�F�
m��N�ҍ���u�"��p6s��l�p �VI%���g�!Y,YJ����<B9���:N|�Zbɺ��cT�Z���{��<c����n��Ԯ�ܰ��ۃM���=ɥi�+��G�:��+߃@܅�Qū|x��:�ɿv7�
�o���t��WbQ�w���1��Ȏy.@��7��
��C��s�XY}�s�%*X�Ό��ϔ�|=�QG�ʿ�V���i>����s�2�'�kOnP���絎�Ǜ��̮��3W����Ѐ���I�5J�����C�"��=:}4��0�N,����=�,�OC`��` ��g�gA5R������!
���7q_����/���7�eZ�e��|�������V?�M��Wݹ���X[��Z�c�0�E(V;e���JQ|;^�=��,�&}5DSŉ�+-��@���p�QM�X���Ը�h
���?���Y������'C��P{.K^ L���r��XꅿHۖ����f�h�yB�� �� �뒿Gӭ�D�%�6U�7 ���>?���,/��;w!�c�Vgl�/�/�_��0�*�����1��D��h��;WΙ�4�d�=�H�CN%���>t�5�Ms��-�M�O��O���<��h��uhjt�"c���K���i��S��l�CQF��Ϸ�Ң�8{�QFPw���ʳ�pr����_�h�j�S��mj�./�Nta׆�����&E=���S�}���W����,wv 
�E>�g����ƹb�T@&#rZ�x�K���;:{��U�����O��Q�P~~�<�$~-j/s�#Nh���^��	#T7'�+SC���l|u�6�B�E�נYB%>��qPޥ�bәJ{��.�rzeJm]v��-���k�<�]���j+a�j@���S
���޼�[j<{�7��""c����xE5�O1�L@��U��{5<b��\}T��U�G�Jf���#���a{,Y�r���ٽ�N����-'��}I��7a�V�r.�>���Ȏj�_��Eu���I�5g�5^�pq���6.<KE��{��g��U�"�9w��Wm^������ -�;� i��
)�ls>1�=v%H�&�;-?O�l�"��)2Q��-'[��9�A@��}�����3C.�οx��"μ�p�a�oP�}ko7�Ƀс��k�|<_�G3� ר�@�F��n�>�윴Z����7�]*���
��Ǎ9��}��g���Tk
���M^�Mz�%x��~m��<�����'y�w�J93�?���f��œ�L�h�RI����<�	���p%���+��&E7�ĭ�8L%���O�f/�N�dO��3є8d=�@���0$����*�$+�b%Jy����u7�<gJ��8K���������vӮ���������`S[7�M�*;�<�Z��9���8R�;�9��$�./����	L��Ëk�J��;�GKǜ�Dy+������qR�D%���9�3����r>+>��9�fE+r&ə!��a#�"�s���46�s��O������?����_��u�����B-�A���A�� p�}|2Aw��`�Q3Ƌi��(an���kĬ���;#ߩ�13�R8���Sktx�Q�G�R���+�}��i��;��g8a�֑Y��T��Q`��.���}�����'jXh�Y���,��3�A�d�o\)sT�e�T�t�*
�<����l�hqp*��+L9v=LRTr4@�ܞ�
nX�</����A���+LG�2h*La���墸|vf���� �"���q�{+�؆荊������F?��_�ÞG��]�ye���l�-�A�K�$h@;h�5h������-_ f�XS�P�6�r^7]Rnk�bbJ PG�ZX]�tb^��p)�ot�䨺O(]:h.e�8=c�ٚϬǹX�mͻ/|G����}�u{QAO��ј94[����o�d� ٢���劫�PsI1gn2ՖG����XN�JP�w��,�a��ѧ��� YV�Kyf"<�m�F��vH'��3�|�q��]H�����z��@���a���J�~�6�?��������z�Bvu��՛��ج�d<`��,�ۼ�����a�p��]���b�M�H�_���B���V�X����V8M�7�C���C�iCf�x�m[�-~$q�(K}�l��'߾�L��.�~�Q26A�wc��P�J(��T��B�b����`6\O���E	]�:I����.�Y�b	*�{�~	i�&�wg��=6/?� ����L�O뼚O
KV��t����Í��H� ��$��$��8q^Y@�.Y��K��%�2�ij�И�@��)/f-g,�G�?	_��ȮW=�kr�6����2?1�2I�N	��UZt%�h>X���X2O�6q{t�/s��:�d�5��}�����YQǨ��`�sXAII�!OԎ���������[��9YXZ�dyr�PG�Q{=7�-!������;�86@�X{���M9|y��@ƽR�xzM}f���jLb�]�ӈ+
�rʆɕ�%�w��5ǂ�i��)_C�)٧�}��ZÝַs�Β�����_OE��Gw^�b���q���\����u(�q~BL�6�j���bک̿�*/2�i���3d9ə��9QX%�oy�@�%,�88�)�Z��d����8aFT��}����3�W<�]�r2����d�U�R�b�.� 8��D(,+6&D��׻D�3��)�2�+DLM�����t�&���s�'�<��ָdr�6WP|�ZVY�G��7�2��جE�%(�q�.:�KJ��T)W3-��񴚪��L�)ϰ<���d
�G�8�Z���袤��Sg�EK�|i×���Ig�"�\c�i�c(�$\�k��t���b���M����w�[xb�gMp')�@oz[���<��~���n�-�E�g�zC���V�K�M����|(p���!ĸ���븸�h��ã���~��_N�-����U��V^�^��Y���J&�p�Ê�5���s��Y���g��|��o��J}*�eש@�������}b'�:
��!���O?m�.I�b�=t��v�儁Z��q��m�����,�}�̫l�K؆��[\�߱i�04�"���&Wi ^�^m��G�KjBߌ -#����wD7vΘ;�����ɑ�eC�=-q-(P�uF"��mŽUh}��Y8ЄJ�j���</I9��(3X}�{#��?�����b;���r������nnz��N}�ĝ7m:�qE��$���(���Gb_�9�1Y�4�`��>����[��6t�$6ǨZ%o������-x5>4�d������Ƣ���kU� ^��+�	N+�A�Z'EMy�P?��Y�p�XT:A��4�Ǵ��ؙ�V�C	��t�^	��|��
&F7�Xb��J��v����m�L��ǥ������C����NFi�z�jsz[��$�m���l�ǁ~� V2�4+{��cN��#��r�a�f313W�K�-�o\�w�4��J\����~���/ �gq����V�����'HB� j,��K�"δD��\B�vh�{Tz�����'N=��(�a�z��A�-�)�"���F�NsY����>�'f�����jey��X�e�#��
0gꔴ�tD�3�Z��>jEw7�h|�<w�S��H��Y��C���I2
���g�G�V���śؑQ���4թl������L69�a�J2��T�/G��.�Q�,Ԣ��T�<{j�wiߵ�^�_L?>I�#�;�ĝ��G�]H\YuL$��8!��U(%������ޙ�}ܔ�"��S�c�O���Ң	"���Gs?%rf�d	����;P ZR�礑���{2�-H]sqKq��z��B���ҭ�L�U�9O�2��U]�IƂ��ݸ׮�qM�S_��V�reXeg�w:+f�e������M1tyF1����&m�x��1��nh���=�.;ԯ:+�[�^��kI�.��n��$�"K-����7ۃ���Q�L{+��޶�+�`��y;�%R�M��ɲ���o��$Y�)�٨v�;?�M�a���u�Vu�[���*	l���b(S��y���o���T*�k〸_�b��3yx���N��M����M9O�����ܨ���Q�fu--ǥ-�H���(����>k�Pe;ΐ	�^S�U_y�c;5c�~�B��1TEeC���Es��E|I�I��߁�^�Q~!sl͗�Ჷ�J���jC+?�����ߞ���^F����?O>}zΥ�Rs�$��w�̓V":�Hw���ɮ���B��xJ�Qt�R�dLW/�"�>爷_����V�_�*�V��hO�4L�z n��C�J]b��I� ���C#dˊN��5P�*��������{��{q.�y�UUU�&��v7@ᇛ9nb��[ 	��C:}���Y}Pqqq��l���k��ví����[��ӯ�B���<�*᫕��]�&����0e��(
�l�`:���C��]����+�yK:�����	ZL�fa��so����;���@�����`���3��:Q,9�2s�Wc@U�OQk׀��=
9�!��`H���D��)zza���_�^FT2�=�����Nae��s�^�k��;�_�n���#�ys>#""�6�%��S�[Vݳ^tyq���Iۣ�ݲ��Ǜf�n/G���~�T��X;9�8`#�PG��9�{1�+`��� -5F��/| f������ �3��n�C���,ցl:��/��C���VT�/$�|��4�`6�-�zC�d�b��eW��N}�/D�E�%�8vܛor?�u��|��� �C䒵�Fl���(�H��g��V+�o�c�1���E�k��L�]�;�$_y�'D~�1;�{<T2+�uӛշ׀��s�A
N����Pf�80K}�	�%�,zk�7������~a�:�g��u�7m���]�o:��Ye�܈t�a��b�i���������[nZ��~k��pR��GGG���si���Ph�����5p�K_�KRV?aj�%�����E&��%&=KL/g�'e�1,����B�;�H�&%��q1/}�30�w<��9�;�,+k1<{*H�oo�ME>���ʡ�\��'�q=P�H�n�`���Y0)���P��bMX��V������yr����oK?�~\��x"��������g�e��O\���ULN�辭#��p��3>;�jطͬQo���H�B�{d��K�<�d�c������֬���|l5t!�yw��~S�_FN.N*TVQ�>�F�@/�t��u��ee�mP�?q���jS�;�(nV�=/G�r4�A��`.U�}�u/z��ZK�L�`�M,Ը�g�5e,G�;e��+�6�������i�e��>c�X�� G}4���W1���,�gƯ��eT��j�}����v���P#g����z���ӽ- /p�x� �����0ә�3-X������=�CsPfN�����n�@�c`�D=��	(�T�u��Qt�E7SGtعL����W�EqR9��J�P�̑ 
������n����e�5DU�:V�w�W�-��P�-*#T,�Ý	�}ʭ[�0߼���R~Z�PA���M �D�zS��7���/�T���������7Pc:o�"z��m�iΤ�U8���!6�Z+k��-��Ҋ�2a3[�(�+�d=�V��_y�^��p�*k�|�g�q�:�WK&u�����u��d�M^ű���}<�/��;J�5��P4j-5�t���˽_�F��-��
�oa:V�5OҜ:�s�EF ��ik���`���*W��x�٨��M�P��S�U�sc��騊�u���0yccÂ��?Sm�+ϑ��Q��s����� |g��D�v�nY2¨�Ӣf��N�ܹ��wG��`tP�w�����7�Ƌ^���Q�:��P<��((��TFR���ȯ�$kڏ ��[�E� ��U�'GXDq����{%���JԖ	�7�&���XO_��b<g���_�C5��V/lM�ӱ��m� ��5c$8C�_����=�]+�-d=�9rh�l��Y��hB���}��! U��{��?�"N��\�a��u��E^BBI��0� ?�&z�pG�2�`���GI(r/C��`
��J����*�͑�h ��Zd��{O�����1?y_�<�^�]�T<�r%)/�p���rR�sU��|t̟�?J���iQ�<���X���a��]p��H���KV�KfP��޸�R�ʽ3m�' �e����;�o7�+�؄nc��?��W�����<��뉜��x�16�����֌Z9K%n�YHC|q�Ѵ]�"X��MQ3��F�L5�I�[��h�K��n]�3�}��hX}*�u߄yI�D���.p_|�����ůh�{c����}}}��~���aN����d8���Z����u��
�?F;��D��"�~�^f�Q0�v|Ȃ���*"(1���[k��Q5�K0k�=P?�&[�� ��Eq��?�����<��`8z�ja�lˣ�D^̞
�(�bjM�
U)y֞+�Z�$�+77���x=h�N�O)yz72[�wz�ӊ�.�*(����L� �Gé������B��D�B�^C�OΗ��x��ʀi�(U����gq���2%�U�d�eol��ݥ���P�\)+'j-_�J��cyy91dg
zT-�6ؼ�����3�\�����%&&j�'<>�����[�dE��&9���N+��� .�1�^Y�u�~�|ɞ�����=���!�=�������Ya)׍�z��;s�|$A�^��x��&s/�@S�j�8OQ 0�[��<Y��Xe��j�M.����X7OOD��o˻2�lh5�c~�}73��^���)������Td���K�����O/��x��p��/hs�����ze�$ľ���md�g���]:/�\���>)"pez��}84ד���������Hbg8y!��7,l����0�y={f[�+3�����D��&��"1���~��^���I[cn��̻	�C��Z�b���>Y�������E�� ئ������B��ָzyn��G��9�$ur���,�ǣ߱�${�n�9�'H&?��X�g?$q�.�w=�_Ԧ��.�rmyV�|/Gʲ�x�`6��~���Փ�������<��rW-dan�}�H�r���V��d{'�n/{�5�Izd"ܾ��2���wŊ�B��4�#�h��axx�m~aA{{��`b���3�-�<�����rԂ�ۥ\G��@��?�A�۟�n�l��r�궶��3'�]$��#��U��tj8pq���%qO��H��Wջ[ېm�*x���^�HH\q��B�)m�:��gf;Xoo�b���M.�v�=�݄딖�������2��=p���y���pH␿�e	p�8�WXJ��ࠈ4u������a7y�q*��<�`��R۰����ܷ��t�$�ՁC��5'G����ۖ�)��Fa�Kڴ��R�os�uB��-���߅2Q09�����R�gnn��R'��L��J���֫�A�Y��K�&-�&�Vn�gt,?y�"�(�y��\�g�ռ�IlOCK"���6?�P.|����;$�W�ە��<5Vj����K�U������rS��㹴9c^7�G�������J"Oc���O���NΌ7�L^��)�����4R�Dn;�\#�˕�R賣�$+%lv�����X�=P͛�P��+i"��j��5߀s�/���=M7�"��7_N������;1HG�}���Ҿ6+F'cAd��$a�R��Y\��2�}���'���9�S"ǿ@Ù1�(����5R��s"�ڌ�o7�Y,��B|e
�+D��]�����x����=]��㤥��Ŭ�� ��˲�_�&߃jt��8�X"�f�Qo��H�Ym�7���5QY���^��H�+���43AZW�Hrl�
|�].|r��1K�S�Ҡk�_"����"&T���G� �����|fh�VQa�րx�y��PrgG��4^|�C�����ګ��2��������t|����"us.��>����x�O0z=�?����i��aۖ����s��&~�B��Ҝ�ZXE6D�FI�jV�:n���hL܎"��^��'� �%�"VC;.�tt	"J_�=+L3�j][�� ������_��d�Y�jw�|h٧��iS��Ze"�!�e��pp+��t�|�R@�ݛr�o�xV|��'�,J�b��4�{	���Aɕ<��������+�  �O�3O��᭧���ԼY=қy��� ���'�]�9���N��nz��Z�f�7���+�kVX����Pq���UT�-h��#�A��;;3	G(GJ���#�u83��W���}q}�Z8��?&�#�0�RC��N�P�r}�d��aÙy�h(`��ʵq���p��PZ�� �$ld���zv�}�1%�(Q�p}�/D�=��8U���"9*��.�����y�ߜ���%�m���t�F\�q~A�zي��${(��t=�\��<�Ǿ��?��F��1B.��\L��(z
�,��W2r�Y�OT�p�Pr����Ju�2�J����F�N��d2<�O��8����[O�$���JiTXV:�;HB�Cm�d����n�Q�F���Q6وG��&�`�ދt!�\�ܺh䞹v�ۮ�=���^'�.ҕk_����Z��:?��ftf{��s���=r����$}����Gh��k����{�93L��o��떇��şC��U�a���W=<�G��*n�W�0���+k���0*����(�+�@�ZÝ�zj(Й@�Q����W��+*�ƅ�#p�����X�����{%����b��f�^c��k7�������,6�=����ɂ��ŻS����ʏ�_ҾLw�c�~��u�F�#'ve�/p�mGڐ��N�,��:6]�.�#~���oul5�fK�|7���~��5�Y�p��i�`�7��`;b�A���#�v�&k�����B.��R�(O����]N!����i�́f���0�N������`���pM�yj5��vHyYҕ���R�z�U���Vu��N�;�dd�t��2���?�3���Υ�vh�B'��Υ���/����(g�.y7�&߄�61��=X�5�|�T���p/��ņ�lmj)H�0K�b����QFNO,H�3�=�!�\Ts�"�gۓ���r��fo�l���"�_(�c��4y��W/d
'���'H��t�민=Gj.�	�֓��;W�E�)��R���'ٰC�p���p�F����q�2O���_�g-B]���Bm�5/B����G)�����y�#��[�'p�����.]�1�����<�Nu���7d�\�5l��SA`�R���e�P�z�[����2�~!Jn~�o��T��H����?�� fr��R�d>�,]8 �&`���>�Ņ�[�6� 7�t|
��ŎO�π�f�D˪`K��?@���g�%���sҮ��,R�����Uj���cԓ��a��Z�=�N�ng���;? ��m(���E}��.P�U�ZX�b+Υ2ǂ,TG�&I��a���	�>f�M�f=������hL�=��H^�O���r��0��Ay��D��w��J�Z��������mR������*��d;�|�K���L��P,)�N����]b��.Dk��zWfS�E��*l��&k&%�<όeG�ޛ�]:���)����n�kiH��-b�SQb�L"��2���y�G��B�=�)GK��/|�2���	�N���p��Y�)�iЊ*q�E��R����X���`����ڜ��X�oGA��L!�OO7����І0d2��>|9?2�ǟ�-���Ȋߦ0����S#�@Y���Ծ�?�78�nB�7;RNcd��ހg��Ԯ� 15I��qi\����o]� '	�n�+�P�nFя�78Č���sH���1A��
���N��??�:A�3����Nhw�̶f�Y�]�F#-�G���sz�u��g���\�單��.�������Ԍܐ�T�x�m�Ō�g��u?w��-���'�����3��\�_�=F.l
慠���͚��ì%o+4΁�oӴ֢�V(¨����*�ѧ5wj��+5}w�Ìnx�w�Z4\����6q�,�P#�Cы�X�^{�jn�Gd�,˃�u�j�������8v��OB��fv��s�P�6(	<7�(��+���+�S�{��Ət����K���6@�4Z �B��V1�.\njn�O�~�6�$�ZB��,�����I��_۶���&�R�G)h?=���9�Io�!`���������隷�N�k����!�^�;IX�:w�Ëul��<����R2q��E˱ų-]��ϐ�$\i5D=��;�巈����:������P�?�6�}��@Ģ5��V�B_��0��(@�I�cg�Y����)(s���B;C�A<ɖE� @�%&>�ʼ���;�Ve�Guy���2�ZP
w�ۺ��w�kޭ�5��֢t��̶�b8���m�K���0�P�m�pG �y�������R;1��7���6�)!��?�����F������?MU�xFڕ�*a�݄�,i�>$��z�!����0�2��G����xKq�P�Ҧ|��Gi������`����V��ԗ]%��C߻Z�Mǣ��HobH?�Gh>�ta؂Z��!s�[������q�uwgM�2����.�_� FIK��p SGR�Y?��p#��t@Ѱ`��慧*c(����b�r��T`�WA@�\��{�S�O�M�~�i���	�[�X������Ӟ��T'v����[�r'׾�r볿��N��HQ[8�}�-Qp�ݥ�j���\uU��7~o�����'�6B@:�>�BS��>���J��4񇗾��T���J`	l���]�K����T�7���T-εĝ������j�����5Tl��r���7��(��?���2R�豌����$yC��{�#s�X�hN���iέ �7�
���F4����4�����.��skYt=�����N�!��.z��c�7|$��4�,~:Xx��s{�{W^"p�72��滿�nՇ.����ٴ�)xt�%B�!��S�����304�P?P���6���>�w���C�nr���>?��m_u���9�k�2t��������<�1�A��%!�7�B�&��%)�k����<�y�@U��Y.��q�I�ʜpaI�ӵq�5�X.�Z����.��BL����f�n��^�bY��'�az����j�Ԓ!�n@�s�x�s�On�{o�F���I�.��w�ځE��͡p1o��+��$��:GR��7��r6R\!����4mFv�r���*�m2�ܙ|E����K������h��sf]C�a�P\!�Dq`f2�g�;��gD��.̙�.k����*n<�c�m{��~�M_�bn��A�w���c &�<��3�!�|oz��zջo�&�,8F�R/���C�vo&q���k�����l�z\*Q�F��������OJ7��5p�N��>��>��o���X�툾��,t�̡b�Lui@��st�5:�[Ħ(�u;8�ff�j濣�_#��Q�HYŕ���k4r�h����|0�]���yX/�׼3�ļ��v�mLwhy���䐏!���./T���|����/X�@t�SG�Q�Jd��/����햺л )i(�o1^��A�d���A|������`�_3����d����Gtvk���q׬��mm�	[��e�,��)\��Ӱ������O�1{���' �
d݉�^0+��޴ ��]��b�^J�E��K�W��|W�w���r��G���i�O��}J�P���1��̮ d��W��"6�>H��Ƶ��������VE�&�:�s#�
U[w�sc-�P�C���xZ�9yT_�(��Tq(�,os���'�!Nii��:�����=TA�w|�Kؿ,bn�]�*�7��	9�P����b������Y�P����ㆬY1.	
J#����%&<�~E%좜}�H���� �{���N=L�_mΫ�j�wmQ��<����*{�AO���Xk�*Z-Yn�4:_�e��53@��˵m����~Q;�u�Kv�����3���̍ v}�63X{�=5���Xص��ؓ'��r�ۄB �D� �(�$y�g&�����U������i�_t{�%��NSc�	��b`�'�I �U�n�?��=����k��q
r��Z0Q�v1��h��V���M�i������5;t�X0���u��f�s���ʍ�b�Ep7�*�UW)�VWi�!�%�:}?��׏�����/�^�X
X�wi��_7�"����2�
��HUl��݊p;�\<���@��l�pU����.$�Kn�����������������ӑ Ɋ�-���:Q�_�։�xy�g9��lhM]p��
����s�(���-v���X��V���΃���[Ý�x������y2Èc���>�:������8�n;>�ـ��%eL`��B��B����������|��ܯ�_���3����f��Q��]��Z��3:�N���� ��Y�c0F���p�(�A����
B�S/uE��q��*���R0�PZ�#(<LQ���R	K �����1�d�X?�Z�rz�\�&Z�t�=�� �K��թv �6�+�7�P�� ��o���)�xr��R��(�d �ʙ������q>�O�֨{��n�$��Y��������*W!��$>�ɗ����T[��91���}d^��QY[�].co3�27|��G�yF��bA|� �m-�K䖕c��~�����#9f�ѯ�[V��z�MF�R�T����4�0H�S!��	��!�p���/�r��\Ph��j�<�cI+tfF�'�ͥ37.�n,�|?mz�cm�;K\�A�����tC�t���@ �}]aV��g�LN���{w��bak~���fe^�]x&�C� �5��l�ξ\�y�1�����5�Z P����=l�km64����!MV��3�qnE��]������u���m��#ٹ��ݳ��R��|�.�����U/���	��3=�^��ҥ��8po�$��OX���F�����{�n����8�|h���Ջ�2���1677�tb-������l�Vn�sK�˅Ϻ9��8�^�N_$[�ʌ=*p���g\F۳;+����

Q].Ժ0���2!�	�W�{އ������@�V�p�&�O�4md���)F�=��n�jV�(�0���Fwwu����|�?�)��<9�*���G�L��1HX��l\��I#�n\��gT�G��8.n�9�0�k��Uv]KaI#h`�?ք��y�휺:;Oʖ��������׆ۇ`�_�%*UZ��x q[h����@��:62O�3������2R����WKKK��</2��k]�y�1�1df/�g�-��Lv�
�|�c����cX蹥�@P��%Q����c(�lη�u��1����[���/�v}j�e��ua�z�d�w���� ݜ�u�9��AlB�x6�gp'�6�L��ͫ����z<�k�nX�m?V
�q����̓XZ�.)��Ar�O���w��=�30|2}ɇ��� ;��<3(�N0�H��ȈO��i �\�?\o%��aW�P��T[�'b�[��	��d*�C����2�ak�|�Wywg%��Aaa��mP�~��bS�f����K#���ocG����
\����PPX0��Q]gW|�J���V�M�8���|�i��<"���L�������0 
vj�qp���Vv�q/�V��4��Z�����dL�WE�Qֺ�� $�"��D���Y����	�-���%�fM����hX��m5�zߩ�!ߏ����p5�`7;Ȏ�o��&&&�:��/�ި���Q���Qi��r�n����C��~ܭ��=	���7��?O�=�p�s^�{��V`3&Rm����� ���vpv	/���z��7��z��*s�o>H�"���6o|��L�׾����0�̛�����Yv?xW�Q�n��z��|�����m��ӇH���,5��b�����5�<1�.�ڭ�i���!pT�D���/����Bd�����
��~��po�W�5֝�y!��wX�,�0	�΋�k�%O�͟��kg��>��g�P������g���x툥�*�B�s�`��}İX>����������4y�Ϩq�'Ɉ�E�Zjjo�i��c��O�C�Ǘ�F�{����4t�����ׯ'���c�/�<L���n����U�<L�~��')�ia�n��X)���s�|�`�����سѧH��F�g:�=�k��6���]��q�y�� ����\�*����T�A�ʅ$x)u����{��C%�#�������L����-ł�By��j8�K^�7�{,uֲ����Y$�I�9J�B���w[j�<������R[���w$Գ�r~	i5lΉ�@��>��G(w!�Z7�4H��U-���1��{y�#�ý�բ {!P�Μ^+�zV𕊡�P�uǣ�O6�.Ku��#����X����L�A\��wZ3�����&
Q�V���k�+��mHx��qWf4b�Ap�X7��`:�X�q�>Ȩ�"VX�I$�z�۵�*rz��Z����oP�!����T��" �Q>	\�xR}=�o�vlp)��lW0>�K<i�V��~��[�^��`�[xM����C�����JE�)�Yf��
�뤞8��4�K���!��҅��U�)B������8��b����l@,�\�ű�����qmB}��=�W)#j�N����B���4���]�����ݒ����-Y�G	�'{�f���i�vw�[�\�ᓵ���
��gFЅ�����t�r��e�(��:q&���IM�l���[(�VރusR��1�u\?N�/�C�FMAKㇵ��N'׀ȸ�\��n��n�Q��%��`1;�I�lf�9r��;Ǉ��q]��3D�?¬��TTN[Y�9^��
eꂠs���Xc�A�� ���`B��.,�7:�w��Oǭ�,4Lk�h6a ��7�J�̪>J���$z��l���-�gD����q�e�0���f�4w�f��9_j���M�����q�7 ��FkA��&�${:7y_�o�7���?P����H/TL�vR;G�s��*U�˵�	����Y��.b�\w���oRF!'�Z6�z��X-�Q7��� �h^��1<l�EDK1��;/����
z������2��ߵ�8�y] ���������t�Q��I�aGH�s~�Ƒß%wk:�����K����/��Zb���ȍ�
�Ф��s)�^��-�i�A�^֊rU>�%g�3�<�fXK�X��������%%�����%$������f)�����
��o����Ԫ�llm�H{�L��?)���a�M����Z����n������{�ԹM�x�w�Z���/�������ź�q��f$�Jg
���R�� ���􏷌2�1s���v�C�"Q���'5G���E��(U��o�w�j�ϸ:����]\�B:)��?��̸��v5I%h��&��Y��n�cG� W�_��S'�|���+���P>�뭂0!���w��{Q��7�ߒ���5uu��O&��˒�8�w8�kk½��)Z�qN�KD`Y�7���`Y�S�P��d8�����)�̌K�#/�J�ɜ�Xpӄ��#[W�_��Ȥp�a�e���'�l8V�n$4i[��ihv�r�]I͝�W�.�;6�X+P�"�h��("'�����qPq�)�rE���K��1P�G�7r��(���ԫu�y��L~�I'5��n��28[ڪbr���iӪ�l!m,�u����Ů)��x�˱1p�skk+�?l���2�y#$�o�GiƮvY>�{�{^1�@���WA������YiPv�sTib_�V�io��O�+��V��f�Pc�����^w�͒�g�<$���=��hr
UL�1���	X?�͙ܰ�5�49t���Q��,④-��ߣnl7-�khc������NO6B������s;�2���7bV�����A�l¶}�S�iõ#�X�KN���K�a���!�=m��*���6��666��LZ��<8������i��z~���[�K��@�iM(G�9B�&'�N�Bm�x9^$~�޺?d{<�(�{���p�AG�<���V���^i�K U����;�{�ԛ"F	3��v�Rd���dtC҈.���:\��<��9��@�XRSh$��+��Н�U�a�a��ߩ����Ӭ�C��n�@��'��I{�������Ĭx�ez�Ԉcc��lVd�ovk	�\r����)��F�R�	h���G�X��X`��W!�o���9��	�j0�8�<"�dZ�yH�����Y9ۙ�R�`:.S�g���>���r��>F��v�E��W_���	OͺP��V8�8!3�:j���Y�3]�Q)}��{4IZ�8��'Ú�$�?���FT�� ���>��/^X��?�ߩ.�߻+�؏:�~�Ց'W��8�q�l��O�.;�;4{ď�z[rhba�9�Z*���kCw�4���b]�xHܦje0S_m�YC��Y��r*<�U\���]��ΫV�#���6�f��x�;b�i��P�c�ϊ��˫���M��(��y�XAҪ�F䇣ø��w�:��W.N��<���}{��8o4e�V�'�1ʹ��=��B�m�mz&�"���+����W�����PO���3ܵvN͔�b3.̓-�ܻPC03mj���bj��Me��.�d{p��6?OE;/'�$���P�b(��mk�$�X���1���L��]�d�yw_�&�%��T>��xU�Q�Cޣ���}^��e5Μ�k��d���R�qԊ'~=EA�VB��RZ|X�ہ`8@!'@lU�H�o���m��_y[��-n%���<AY������9�U��g�;���oi��1v��+����qK(�r�=���7YL���:��uw��c�W���P:��H��s�ڡuW��|��1���ϒY�^�3���J�׉E�R�{W��U�~%���q"�	'�ui���/�\b�C:����w�J��|�?�����pf��x���?A���b�����Ny����9an����ܨwjhd����G�lش����D�=򳳳aYӆ��lؕ���x�~ M�O��N��l:�j`��l���U����%@0��s<��.����y ��[ya��3[!S�e��Ѝ�;����ף��hN��|k�/�OH�xR�����g9�S׹���U5��g�>;H�Z{�L�:ֱ	���]k�<w-N'��+!�N�r<i���}[���g�L�Y�߰�of�9:���LL�p�Ȓք���þ����n�?�Wđo`��q����.a�Y�{�����N�W�+'�S7��֠b�~���@������j��Y�B�)zݝ�?[p��h���>�	r����]��Y�Iςƴhz�)��V�N�R�"O�<�Q蝀bQL�Y�bS�k�ӯNr�ӌ���͌
+�Y��U�����X�[��6�鍐#�k�_aF�ŋG?�j�!��`k̊?GF����n��#I�K㰩JVa��3}��5=�,��̍kߤwO�<LN9��U�i����[��x�L�x�9o�����'����W�9�~�'�nZ�6M`���R��F9=g"u��Y��f����K<xF]�u�:������AB��Վ�}
LLM{��*ӎow�۝gs8�;;m�o�M��u�졃�M�l��%��;W�Ks\����b�bi���gT��7��bC����HqF�CA�T����(�C�P" DD:$"%"MB ���'8���~|�}ǥ+p�����}���<������s�Nj>�*8��c� 'r��*��ϥ�	s	B��+��]~yb�����(��/9��f�����*���?���7�f����<a�a�{]�!��:�1Z�M!׷�qf��%S노Yfh�5����y�!���h鉆�u�zN�)x�@�T^�Q�t�FY�܍xA��qͯ�����"��=�lo��{�`oΪDcŪ��j�d���>ʬ��+��ѷ�G�.�֔���96q<�*�!���)��njBO�V"�Q-��L6�"Ï*��z���+��5��P��{��~^=[�tRk��5/��P�|������v�f�D��L���X��_uW[)���f�����[r��`�O�b*�EC����SέԸ��k.�|�,�OLM�Np]�o6�\��Vޡ�2�y�d_s����;[SQ�>�M������ֽ@�#���r%���hj���FW�x���C0���^}�	��p��˂��ƶ_ŵ��q�ŇV�既[>�ӖN,$�V�=bj��>�����3*����Y��I톦��p����yIt�҂o�}�m�X�$�\������ ��|���[�+IH2`D�!���u�	Rl��￫1��a��ײ&�S�a�Y����+Y�X��g��'�������dRc3<,�0�}73,���9��pDB�bE��>MI�I���Jz0,�޲���;���D��h]�����:�"e��i�����5�8�m3��cB��O[�F���g�2�,����$����)�����b�9K�baW;��N�\�o��P����":�ͩ�Q�Sc���gY�m��?�C��a�YHd々�w�@�i�������S��MX����*܏�u���%���F�x<�P>۩Э�OOO]O����F|~3�v6�؇�a��������.������_+�իB2��E^~��3N��%��^6��l�#��:�Z��L�����l�]���T��*~q����NT[Qp�&q7�v�a!��9�$�A������6λ�Uv�Fъ\=��o=,��� S7�{�[:�E<H�R��ϭ�x�P�%�ݞ:M�匏
���iv�:��#8"�y����6<4
��8�9��_�/��獒ڒ=�O������.8IK۫ɴ�e@]e�o�>(�]V���D
�V�te�A����GYͫo���L�]tM���\ɭ�tU�K�;���?䳯4����P�vL���Fe��e[��z��e��G��o������M�۳j\�v(���q9��[�1�������]���T�!�L���'��PL��E���ô1rs����P��yX���U
�mM�Uǚ�b��!K�
��(Y��f�t���M��I<���r0Ly8m�@�ǌ;��Nd�H�9�&�ɛ?�z���
�������)��0ٷB�J�$Y~���HLBF�hK��n{]��G��(l�ХЯ����g��^<I���H��{C�(|�='�{Ź�zO/��@����<�xhvMU�����e2SjS@���L����K��;��6Q�g��ͺRU���U��O8��[u�>|�$BAn�A�uaSŀ����v5�K_�j-vEχj�b~����а1�zeԥ�#���iWVծ���/���^u9�J��*eveW�;7�V��+[ԇ��~Fh?�?�!ʩ6�g���x��A�Q�?����<\����z�i�s��.g(����Ѩo��Yʪ�����`y�٨Q�� �n5;=}9��V�獋��o��2��t�/P]���)�ei@e�tf���4󲳋"Jӎ���C��=��V��CD���r�g���و�s4M����a*2�s5�U�%j!���W5�ZX�\i�4���W�z�',������&�#{���7�q�^}��n;ƿ�}K��Ȫq�&�d{꬗d��ʇG�{l�|X�T���Fը�������u�3z�G1@���m��8��Ol�@b�3/_�&�!�.]�F�G���8��FR�y/��A�<�"�`���� # �hML%��Q�q�괻����!�oY���z`��!�"����w,����:����h�lx&��x5��憃hXF��_����j�Un�>ut���v�[���T�(��ɕ����twi�����!��D�:�;r���p�Q�5�<$��a�Z_�m�Q�fl���Z��]n;JU0��F���a"Aa������+L��
�U�U��mI�F�VЌ!��2��F#��u'ֿ��*3�֣������u7�fBO�1Uo)t�k��S�3��!���SEc~p��me�Usu ����Bв�i[^*'Ղ�\������R}jd����U�g����SU�TZҒ2�HzMQ�ow<��2:�]��
+�8�I&��EE�o��6ځ9���㸌��Af����5��\�`�ѱ��Ͷ򢛩�G�p,���������|��I'�D�X �����(z)�c�l{�!�����ݷ�!G�{D�{��vu����JxwT�n�J.�S���$(��+��6,��S0��.�JZ	�/ӂ3��dCŚ���Їڙ�6���I�P6��_�JVj@9ЩQ'��P����.Ӕ�]�_���z9���[N���k�����lD��{��سh	ƥ��k�5V����6��ҫK��7��v�+PmW5���qb�L#��� ��,>���˵�b�(]��T�N&�u(��d�H��AT>oxA=S�C�o�������Y�<5[@��>�=�����$pWQ4֢��)���ˌ!c(&ʧϽn	hQ��/X�*yx���e��܀���uI����O�o�ꉏ{e�þ�TI��_(#��h�S�C	�Oø��c���p�?�1������0R�\c'q�0��o�=��H^�d�V&�y��#���v�Cy���S���;�"~�}|�Y��l>C�tDa����%w�E���P�b�VWkᴛ�\�1���l���q�U��Z��`B$hF�G��&
�U�}��q	�nj���U���Q
��]��u��Vt�W�-����,9}Ɨ�b��z��u5G,l5�y��ai>BF�Ү�%d�T8� �̀s�zM�=�ݳ����|���S֮V�4�w�Uc��V.#����Q;��c����L�g��� �� �ًN��B��{ZT�����룯��������w_5��"�n~\7?�b�6�;�v ��Z�!l������SU$!r�%���s����z[:?W�i�i����؜7�I��F�,��޶��đŕ��8T ߹�ӁWm�q�v�H��'�P�`�a#�YS��_�"L���Qg��da�
�]�{\_�%���.:��T����>��� ���,��k��I���%z��6�sXͧ#�/B���V��T?0�A���F�w�Ե����G4���tm����qM��4�J&o�y=E/�T��>�rzF�[���E$�s�@��'��u�������Q����L��M��ٜ�ft�j��0�a2%!9��c�5���CL���˟�E��8�3���=@{s���:�vg5�u;�N�R�ht�䏫�66mw.G��E�p�{p����M�*�\&84�%�;F�GYِF'��>|(MڜFӖl<�.Zgɛ�Ql�89�Mx�M���.E&m�V���j2�CM�x2/b�1IQ�S�=CmduI]|G�O�� OqT���Xdai��H�]�2�0�$X�(�=mccHPQ#�ȑԔۀnb-c�T�
B�Ѫ+�pAp�1�����11�"�{�и��f=�C�����_�l�������J}4��Ғ7vi4{ۆ�h�_^/ ��q���<�eNA<��b�AC��>�Á.�7�CB��:���k���ʘ�5E����-y��/��z�ݥR����Xa�E�V�SU��H�(Tߜ�g*e�5���媌��-S�<4��5��>���1��*9,������1O�0H�꾸ԯ��ts�z%�ܲ�:7Z�4r�wo#Jm���m��^�\�ncC����;��T�~v�A�������v(���Ņ5r��T^�Y��wvE`���Am@:m�PP�S7�U���E	.Y�l�w���λ��M����2K���sUn�8Ӕ\L{�����؄� v�L�c��3�_B�6�`�|���U%�E`���1���&���C���&[����Q�;X�6��O"��j�'N���Ɍ(nS8������Ѿ�d������B�/�¶M|�F$<����k�+���������Y�ɬ�x sYg٣�,�>Y��Ɲ-��qZ��q�3�&�"UjEl��c;\@�O���u_˻hy��t��IY��ˮ��$~Q�����I���OI�კ����"�a������!+-U�l�_$�þd��v�Va(f�B5*�n�Y��l�)�w=V���ܤ��g-o�duyѧ�L?�e�f�z6^��Ы�����f�P��i�C�P�N���E�W>�u�<�4�0��ӯF�UF�,��Pcq�LK7q~=i��m�Ro_b�6=]fr���D�i��5����ι0�37n���kKW³��\;
1y�y�$
卝�+Bu�"6V�M�ٌ�L$l��CH�en�����eX�u��0^����Y��hY��Ш�ML,YKkĕ�@xa`mm��$��)::�.SF���8�b,�\g�����k�/��&,�E�?��ON�MM���D��(��M��/vv�c�b��)$�>"����`a2	�*��T"�1�!�u����x�G!�f���,�>�V;#3ӝ1�I�	�GC#� q Y�Ѵ��'��ߦ5�D�n�$���'�0O���Q@�Ǆ�XXf���k;��k��1�0?[dCÐ���G����鵕�����Y��������;>}����}L>�$!rm�	SE�ye,"���>����4g��O�[�����NOn{���JCC�E�ׂ�����7<Vp/=e��.��G��{}�f�&F,slH�(�M�>T	�;[��]ܝw%\�˕a4VUJ����ƪՕ�ֆ�U-�zK��$ !�p&�?;9�k��X�j��8�����`�I��"k���m��,���i�{W7�W45�0V|�"����T~��\_c�v���rB'����W��Խ0d;1>����UK�(��`}3_�m���K��~_����*���;�)�J�" ;� }�8��3�a��SA�,t����Y])	4~đm?]$11c�qp.��\�u']�����]^LӶ &��1�-��YƥU2��P����yQA(s����CÔ �B�)م�t����FSw��Ą=���5��TNN`�d���X�$$�G!�$U����
7<��n$�_n��ذX��\���][ч˨��t�l��=t�WJ��}���f���߿*��p2?�144|
"��8[Ŋ��g�C�r���ř��d ����UU���	-�T�ǃ�R�h����K�Ǝ5ön���}�Bo~)+/o_�JGQr��&N �dHJZ}|�*�dg�p� 8������ ��c��)�;4B�??YKwtpHXo�ɶ���\�BT�����}c�b�PƝ�������־�$C��{�e�g7;Ɔ�����^��#�di��X ���>!�%�r�Y���W��;�|���~��΅���?ʹW��}�Y�b۵ a�N�d��[�9���LV��ww�����x�u߹�Jj�j]����	�_.����wI��1+��J��x�I@n�Pg�>���_��]w�)f�	ZP�C�� Q�!����u�D�E��P^�Ua�2�mc��� �,|�J=,ִ����(��P��zM.0�N���Ex�X�LV�qi��Ϳ��h���0�	U�V)1�}� <��Q���S�I�+��}I"�E�Xx^}yɱ!خn��11x�������g�lC���l�ا�~����,��&��BV�"�aN���6`�e2�P��ɻ���vu
z�B�	�y׵�XR�����ໟ7~�%��uw��������#���H�G��lI�������g�~��i�vL��d����aZI`R_Li�m5�Bs�KK���T� ��<��x��n�Q�É���fz��5���pA��F�$��SA�K��Dӕ�&+�@�� �p�֔�v�qg|�{�{�Uf�ֵ����O`���7DO{�ͮ�՗I(֕���S��[�c�6gx�U	�'��=FZH������p/@o��s���*�B; 4�ں�I:�Z*�MH6�C>Y(�#\�b�]�ܫ��,�����[.��g[*r�n���d��)[���}yiy����uE zV*��/Q֡k��D���ٔ�qI��Z���o�m|���q�������>���H�G�?�����$�#�<�iA%�Q�^Ĺ;Ӌ���$����5�s�(%��J:��0�@����5��<�{e(%RεL���wЯ�5��[v�_���q{��?(c)?���_�����b�����©���3=+&-YZ�s[[wD�b��v��F=��>����o࿁���o���������_����|���j��r�J�������Ʒl��_i���%�v7, 4� �Ǻ	��O�5�J�ƌ��l��?o��I�)GZ:�U|��6�s\��:�C^���!�߱C��B�"ʎ�������ح>#�A����t�>�O�-���x"�J��a�n�B�`���H�:VD0=�@eb�]����9�HBj>>>���5-��ߝ��u��|*�{O��0읝��ҫPx~a��#̵���EY{_����]���+URR%ԟ�#�*�n�Q8:qWi[��n����¥?�l�Y���TpF��,���}�m|�~{P������Ϯ�l��6ȏ�܉F�������݊ɻ�␰T���Rs�~�o���ˍ����*u��;w�s��^��rb`oM���>!��ig���L;_%�JV~���Tm�p̧߶Hs�A�G��>R��N�x�.�މ^�t����1�t�n�p�H�Z�!ӊ�w_ٻ�f��w@͔���C�QNjn!QV���]A� 3ک��b2��͸N,R8��}�\P����;�e�S�$)˳&���-�~�����ږ����;9�"v7Y�*+0fؘ��CE��~�芁�:WteW�}�15�5��S�P�-vB=����*|HUSs�_�����'(���{u�O�|f���N乢�4pE�]�������W���FKO���{�
8�����2Ok��P��][��{���V"�D�ʍl�{Ev��>W0Y���Y��������ʊPDb6��,�n�kGE�+�#���K����?[����V�����h!_۲:VzG�8u9�ﺞ�Zee`t��Wn ����T�"��T\�</�|t����`����G�?�k�:%=N��yx >Z���c��VNY~��;����-2G'f,���X���&Ik;lv�pv�ܹ	�1��r|k����] 3��Y�>�Un�����H�:���ł�-�=��K���L��k�"�`�te ��حDR�������#�����t�_�mYP)Td����Y��%Y����#��mV.�K�sl�V+O<�!="�j�R �=���׃H��5|���k���Yw����*=��V���JJ���B������������֯�R�94����A�w�V�:��&�4�I�V�԰�[t+��;F�|"�����G6ÿS���o��2��#5����i�1�Z_܂{.ة�b�7&�����5��)��� ]fϜ0ɉ���Z�ۊ���@�9�ƴ�r�)((��޼���MY|Ш~�L�@�a(t�}@_��6�u����0�h,.�vkQ�f��ŵ�Yhk�Y��:5�x�`k�9�
;bٺ�h��+0�U���s��2�*ȃ�W�oxQ	��?��;���|�]�$�P+x�W���p��~��|�{j���I�3Ƶ�N��O먎��oU��=WKR
jB�?�Y��A�]�栶�g�r�^ �6�E�}K���#+�"�����O,Q\͛:!*^c�����$�n��~~�,�=D�+���^6%�h}�����W�ռ�ܕ�u������ˁ���Vm�q�##�����Q5�2n ���H��w[E�4c\R����O�؄��p��^r�ge*�o}}3::Z�u<%�����%�()�Տ������404�䯓:��1�2��4�)��WS�����333�c[}�gtB��ɐ�d.�H��������/U�-�����r&53c�ݔ+�ĶDI���4�Cy{,:���/e�<�1���n����/�*��1_�W��x��(t���3 v��xf�k��6�Ӫ�����؋::�t�Nm�}`|���Ｏ��������z�V�qB=WOML8�J�I�jC�Y-�MǸb5 ��%��0�x�$Q=�L=Ί�#���C�*�_�}�0��<�����dL��S����/���k·n�L���JT�O�/�`'ϔ�*� �A�Иf�[3.7��~�x�}�h$�l�(;[,fUp���:�xݲq�m6^���٪f��PJ����Df�ݱ0���I`�q�gv�>��G(ڗm��!��I#��β�sEɼ��j����;�����C(�7�
���齵�¬a���(��i�r�'2���)�Gi;��ǸNM���xM����ېu�BG���rei�aKANg7~�P�JN���R�\O�ߑW!�yH����^�^�Eh�l��n�I#Bw�3{�x�<����_��ŗE���}3����_�x�e�Ĺ&7��y��K�Hi��R>�k����I}ġ[h$���)�U�6�,*��U��:" ծ���� r��
1��R�n��f���z:�L��zv�b��<�y��ψf��ڟ�����Z�7���P� Z��dȌ��m�w�]�z���Vv�?s�NViҴ�Av�}��!H:N�r:��#w��6���J|cy�	��4)��$zN�60���cp|Z��0�b��?XM�'A�5ǖ��_fr�|ѨKHs4(�G:�yհ\I�D��u�a�$h��'�\S_�p(+�=T�0Ò�Y�^"�1�R��� :js�#�ed��i4�V E�B$xHC�����˺���<3l�u^��I�^�ʾ'L�h{�d����Hq��L��=]��/d畞��?��80��6�XHYN��lN�%T�9���#��+9���t�7�)�ړ��x�<�1[�1��\�{_���t���B�W��腛sN����ՙp
�7�ۓ�"��n &,���Kg��n��l��l����C�b�&utt|w����`X^�&~m�I��˼g����8a��d2��������v��\��O� ��A���)=Y\DRR���_�ۢ�G��0G	܅�Z��9��W������T�������O]��`h�c8��8%���o*·�diRq��Q3��^�Ȭ�ԧO��}�,���5�A�&�V�w׌2���ߓs9�To�l�����{����J�4 ?L�`9��Y�;JS(TL��M�'�5%J`�'���Zj1���N	Ʋ�?Y`��b���'A=�W���4���V��w����i��j�t��v[[H]i,;���Q-�3a�sq}�o�ւo݇,ymO
��_��������"�P)o���}&�b��w9�������M(�r���&y���1��*'� �����|���{ۦ�=Ql���htd�9�N���I���HkSG�ij��Pim��϶�-|��X�1�����Kºwm�Zc|��2�贫4�ރ��Q�E��lג]XD5m�nU�d����A�v�;�5��z"znº �3K����<=f:RU��V|��?�f�������(@8䜉��^������>��+󱷘m7:
� �Q�� z�� �Oe�
����:n;���x��s�w�`��H�ҳ��,�#Os�_H�6�^[|�}!/|�J+�^9 �}���7���wŋM�,�N,*�~I�УxAz�=3/b{�9J6f��ˮ��t���z\���z�XߝG)��+�雡S��_���p4�jY�g�B*�z�CM���Zs/���������m���~RT�U�P�S1���⋇q�hSE��rAs���L��4L��]��e2��44(���h� �<v=�z2��D�ߺ��Zq�j���w���bd-���њ�a��!<��H\�NFⓈ��}0�lOx������Q)J�Ք-h�i����,�:�{*��
g>�_R��V|�Lf��_�S�ӐK�����/�S<U\ÿ5��m���9� ��5�H[�q����������*�n���b��x����n�o�W�G_� ���9�����i�*��V����h�������}��$���)*X��,4�9%q���\z�J���>���gQ�>(�.	�`iN�cg1��Q�h�mm6���.I���@i��G�b���1(�F�♌g���3�H�n��͙f�(��X\\&��˗�u�.noss��v�oz��K�����q�2�3YS�yȾ�eo3s󶁁[NyY���(�}Ĭ[.b��k�1�n�6o�\|u����2U��E�ȝ���	��6�r"V�+3/����Ew�9=f�_�l�hQY�q���z���!T n.�ѭ����Q��Oǚ��\�}���������k55��S#D�xj��aL�Q(;efwy�#S"���e����	�߫�+	n�bvG��,T5��ʟA��k�:~=������#�����)Z��͞z�OQ,o�����Iz��~�I)�1T�F�8*+�����555U]]�LO*�\<����?,vآ������:��d�4�J(6��wa^��q��L�o�"��
�/�;��P���ZAYG�8!4zv�9r�+�(��#��R�Nߑ։���?!"�'���j�������_H	���`��
Լ���>���s=�5���Ūm��gf��Z����ȓ|~,�dJXc
�;{���G���d�݇��uO��c�¶�����q��-��)/k�x��kw�W���<�M(-�}�hK�,`�)d�"��#@7����@F�d���+*���V��hK%+0�������ٵ���1�c�r�"��I�d��H���8�}��Kt�;����7D������M��p�e:T3j�l�AOL�pd�u���Q��b|�H�����x���ʔ�w���Ѣ�i�#��A��>]ktMtǸC�����������323ݼ�v��{j_X�ts���>vH��a羶��2�>ݒj�VZ��C`dT�b����2����.�}�Gm��q#$�Sc��|����E>?�$=NP[�%^�>x���&���5e���_�mic%3�L]�ee���:f?�r�#>�ل�.��$n�r.ELy��%�K?���O��i��"V���DͲ2L��k�cWӁB.������`��m֥�zi�>y8�5\�Ļ~=�4�ɪ����zp��ȇx��HdT��:��5���������;ȡ��$�4��'R`���[8͞�;̥�Ek[)� ��9넒�Nz����}|0�!:}�-��YJ>}.��6|^�Ne��EhP�����\؏6k�N�:�7��3��=��RQ���M����f\�r�ekJ���9��B�N���x��܀�*b�_�=�w�>Z�$�p���rsuU���Yx�W��yҮ,���o�mI��-� d���Ҝ��*?�����$�`��)�ZRN�e�,��듪z��b�^6�(�������mBN.o��0��0�V��䆙	����O��z<���9���܈/�2
��Rv��缊������dy��PNn�T-w�&7~шG�h�YG�ht���-�aq�L��+JNE�n�;.�v�ڔq ��I�$�i.�q~����Tw3]�E_��`��A�'W���J�uB�
.t(&t�ޅf�\e�*�N o�6sG_�p5�n�D%��ѝc[�FЩ��u�sjKS�N`NrH����Q�Uԏ��(��-�=�T�,$���Je��Knhc��)%#��%�J��_�h�n�l�C)���i�\�p����F��`��U�%핷s�Z�m���s��W�	R����66e����*� i�KS�6|�O��,���"6q�?p� ��74m9꺞3U����1���^�Q׃�~#���oz�f��Ē���(?�\fxi�� �3>J=�m��D_�zUfb٤XK}�0nJۨ��-V�G��خ�&9���H�T�}X�諵UI��,t�}�ڹ�!�/@�i;�����O��1��8[��9�0M�#�ӸfB���z��H��z����C�E�wSmK���`F�w��n�:j_
�~^;���)���uh�'�J�Uտ=�<�XF�U�>r`A�A�ʦJn������W���s6�mMhw��J�JM�_E+�S���K�!�k��J��Wi㝭��~�>QHq�a��Mit����׭��[��FNhJh��?�s�t�u9m��+��躓1�i�鍍�Q�3�\9�;�Ŵ7�_���v���sX6��!�n�����"|y�W��N��6N� �f:A%A��:u��螾%�h�N�3*�H��-X����5��A�&�`�lS4�j�����5�gƫ�E0�kƁ?/>�ߚ��O(샇��F���z!\N����v�Ԁ_�xR�X��ڍ�� :����w�s�;'����<4�7�O)�>�=_[\�F��8�,l��;��F��̈kH���C�~��&��:��[�S~�����$h�@_�Ik��N��ޫ��G�1��,�ۀ�;�]�<��/����	4Fp� ��<�mK�9��s��47��H�؍������2���<�Z�	����8����w"#-Q�=`޻����-��!0[���'F!�p~���:��Z,�� �V��r�+�)�W�b���C ���
i^� *7bl�I��<O��P����s�Lk �����^0NƳ�ֽcrϝ<9ڬ��������B�"emv`��<A*���*�J��)��l�ȃ�Kf�����]�7W7����G��6����^rMxh���і&���Щ��T���v2��-��"�֎)X��P�\
��a���8�f���N���7�y�$[�eU����<�&����=���6���amYj@�|��sm%��I!�2�8ϱ����Z���~��Q��4��|^|�p���J��D��TB�Ӎ�����#�]���*K�YL�'����|��$�7�c䢛�n��U~j"�
K��G��A;�?&�Tb��x������W}^ʔ�����9�Z�iag��<<ZU��H��<�� *����jP���G���E@���7Xk���  z� }���%\�����Ĉ���iVR�n�~�E��l�:��D�iB~T��e��[7rA� f�:̥�tz��K? 4�U#���	\�+51_�A�L�D�i�E+�s�0A���7��ՠr��������V&� ��D\X��d.�����x!i?#&�9�TqK�4^0�����x�\H䟊���A�[B��nT�J���9)�v�߬H�����9�^0��Ҫ��1�<.n���Ͼ��t�v��Z&_��X��O��,+">">�rX���+�.��c]7y�9������KK��%$�l!���!���������
W�W�ˣ5\"�@o���� �6]�<N7l�&ǜH����Ŏ�Z]��5�m@V��� �Ooc�]� �+1>c�6 �l��E�V*E��5����'�Ƨ�pD��*��-NX����c���	4�:�ebЭ%A|#�w�MㅐQ�w�V�*H�`r(5�[�!����3���]í�+�PI�;u�sK�Eq�0F���˴�=�F��O����'��&\~�����`Gg�$�j!9�d�%*�>�qENb��Bm��ף���G� ��7��bf؊k#���?�	�Rޯ�k�*^�����.D9h�_z�#ʌ����ۿ���!�BM=�����n��%���7*pK}�W�I��K��6��.���#��࿬b��a;�ͦ�ݮK�' p�Yc�{�S�|5��	2�<��5�5��Ɓ0�=G�;�;��b�1�?C����Z2�oC�.0G������tA�ܨ�F�a�Y�f��g�q�8�LW�*j�� R1Ȃ9�;^�#�N�KDyʿ��4��Y�[/���N��7�>���x~4�x�B���� \a��l����_*E�".���"��L�� ������Tg7[��f�S-N��,s�?����j=34���#%0�Wjka�qF�����fE^P6jm���#	5*��[zG+6�耵e�sцJ2�:�(ԣ7%�P�7��7^�|~5b*ϪDN�!�����9Cz9�G����$EΪG{^G.Ȣ��x.-h�k!ꃋ��0<�'|.6!�	�1���Y��ǾFI+�Ih}��Iͭ/(��/�+:SO������cc�p�� ��>X{9� �W�*��|]�c�Q4�)�r�ް(t���
�+�˄�h� �-l8�G�6O'Ha�B?�7r�������	�{#��I���4���+�Ham��8��rX���~ݭ�\�}�|�F��\mT�`����W4h�������W�ȷP�c�<�Ϫ������_�Y_�)��G#H�[O�A/<o�$�b��m� �	
�:���Srn��'�y|��k{���CIE8�.��s�>JK4�F���݁=�=sF{�}���d��	he���O�������| ��Õ���?����5p�oay�1���&�+*��v��ґ�G�9�ށ�n/&t�<����ف���p:�촘1�q�,�Z���������V�q�?��y������'���o�����C��|u���B��3���-"���Orȕ�xFD��ǩ��?t�����̿'�~�~$��ɿ�_�{h{���������D�ԆoR'N����(-ܚ���^�֖����Ny7�գ��*��&�#bm�`�#�v-�M���\�YrU���A=НM
:�CXrt��I�v![S���d\�W[&��n�h�(���Μ�_MW��t�5 |֞:#Q&�ߺ���t�/��ɱ����멩��Cb}*b���?˅�4_[~k_�[�B�O�qK=U��J�NQC�l
���j��{�h��I���H8���u�ә���*5v��V�������N^H8�e�����G�硇��`EX���[	 дt0�u�`���Q1��q��;/j;H�/��tQ�pt�7�2��U"��|�qq���u���ş�3��=�'�tcM��?l�థt�_b��$	���z6����G�� F��.���^����a�YL8��������[Ǯ� �e�N���8�'1��^�L]��5�1��n�}�Vq8<�:RO�>1����h����`]��(?�5����T4vS����۞d)	oꋘ��c��Қ���9V�5ab�c}��� �t��>fZ_x��гP��i�V��Jf���=|�K��hag��ik���֧[��B)�f(g�9sf��n��99����5�v �@����W��tB��,�=�s�S䁅g3 �T�3S��w�UKh�@�e�3�k���:a�[}%���?o���PK&kj�2�_z��_3���J���CcJv�;!�Gc�,O��UV�Ƒ�@_oɦ,,,�)�mL���UV]?��'.�"z��ؾ��-�����]ϔh�ls���i�x0����Z������K���z��ow{@/*vMzݻw�x�p�wt�d�����]�zW����m�����d��4��d$�D 5�:�m���\�E��[�W�Qׁ'��Ŗ��� .�5����C��b��?�k�O���:k.D�	z��!��Lv�G��O� �J�^p~^^�[�����i	����`�����8��@T��k�g�+
Y�ۃB��%t��^`e�ǜ���$��E������-[�ƹ7g��
C�,`���T���R���:k	�a�=(q}e``�`�h���Cʧ�(���f�]੐u85?��Dz =L�C��kS{z~��ٞ�#@ �l�R���GQ�q�ؼ����̴+�)Vc`�_@�ٔ�Wn�?�m��h�O^��)�!j���3!-��ʰ!�f�윜]� G��=�9��Z�|��?6ѱ�n��Gn���퀕��
T��01ė�ϟQ~m��y�����x�,4�.�"��Q��Q�w(S���\j�������-��2 � G<U��>�zR�v�Zw��j�^�a�k�����B���e>/s��񻏮������9 �y�4���G��]�o^��5���������Bu4�q���ޡ�V[�ſY�@��B��'BYo�(`<��t���dQ��b}����7N�.�y�����Gi��+�}UO��)l?�!�P�/l6���\P�Hҥ��<4����BxZ2BN��)��%L����Ԯ-^�5s4�\�6����5a�B��ފwõE�X,��'3KKK�VI ��v�S� ����ō[���8X?������Q��a���M�(
9ģ -�H9Ao"�R
'n����.�����ǯ8#؜̙F񏐮͗��1@�x�� �r��c�3rUZ=QJt�pi��++~^�����|rO�����/�@�Dֆ =l�(��������,A���N�vh�?�]�7[y�?�������vP31����u��ԥ�����K�<(1�	A��飂VF�1J��U]B	%H�h(�(!u��E�hD��c������9?e����{���gO�
�
�[ R�t�y��dO�J��; ��m@�o�8���Hg��4_ IE�?J�^}���}Kww���'��������=.��n�"�����nld�e0��oa*�ܓ�Vo�����p~<�� |�q��aH8�l�;�!;�7�ۛBrQv���
�?��F�ڀ�� ; m��@C+��`���tl��oF��7y��H�{
��j9EP���-�T�V_&�<U��F�~��n��v ������)�r��C����;�e����
����v��
��'e5 W�h���5���'��ֿ�>�Ӱ����h<�߲ Q ��@hd�'+'gLݡ�䴿���ԛ��J��ؕ���3����gi� (�C��7Qh'���9�y6� 6��Jp)-,;`��q�XG��0\�p�N	|�����C�9<�)�֡��9g$<&j�;*�L&?������`�������. ��P��H�rc��I�pO�_�c��q�U��Θ�����'���@�*��Z�[i�z#	ʇ��g蟑G���V(�o�����'�E%�Ⲭ b����B��-��	��D�k����4��|&��'�aN��;	t�1���y�ح����U�Eb�SWף#&���U��kE.���-��K����y�i"h*�<3��Џ�$�6砡	c (��[=����4~��8/���9��c�r��Њh�4G{�������/�Վ��v'.@������?F����?��M׎=>�]ɞH��-�r{�k34=��z��������L�<�a�0H��L�D?rڹh����}���ӝ�X�,{}xp�T˩Rm���W�	.r� /vB?,ׄiq�M[��x��6�:�5�;v 6��P�^�BZ �,�[�T7���7�t��ҹ�]�eQ-C���91�G���O%%U�U�Re���`�·���z P��7g���?�rɇ�:��?v��A���lZ��#B�y�O�x�b|���0x핆�Nk���T��JQYl^��;�.P�/�����67�G�$6����*?���{:??��I��D1��s8ԁ�I�7j�y�F[�.�!���6�����p�ŤL��B�ѵ�5�-%&��{ʼ�_�$��*t�U�^��L�*(laS�8.5;a�4k���d��9ӭ�z7���\�W�p���(�}�3&�p9�U4:��ѭ�fd�;���hu�U��9�؊����f�4F�B�]�Vow8()�!�S���A��@��n)Ơ���b>��zlհ�|��JZ@��x�'%�*�mGC�Y��[ ��y�[�/���� �����#�A7�L�5��Y����� �Z���6MY��T(/x��z�d�Q��O���z|��+����U�&Z?��v)H/�Ӏ��T�D9���j !"�wֱ�[��%��S.��l�-x^�kV�����iHo�x��R�>h�������(�B6���)7��zm{ (�ޤ`R���qlR*2Հ�������N� z��Z3<�L8D��a��{#�}�Mq�TC�M��߽tB�s�>l��.���xnB ���?o���x�+l�6����� #!�5�یګ-���5��@>��ݱ������W��hc�|�D��N�*h*0�w���`��/�zi/p�$D4� �g�i��+�]�HCS��P���|��a�	�3�f��K��~���kGd-�z\�-� W��t� 7� ��T����A�A�� (�ƕ7˸CőР���>y+c�NEI�����8�k��� �-;0k���=V�]c���m>�A��f܈��}�z�m�{�`�f��e��z��#���<R�D$�%=�|���.s�3� ����v#=�;b�U嚚�0�9�BS�v�D��p�i9�S���pB��!5~w��i�
@���~�8 �����$�#Q����R[��-��[�3���7�$[X{Zbutxǁg���P���iQ��E��z�GN�k��v8�~�x�ݶsB#0�#�P��I�Cb�4�Ѫ@�����@�R�كp%�W��0E=0����a��@ի=����7��ſ�W��Y���"tU.�G����Q�G�)/���cr�͒p�6�0�F!ٗ��D�DRM�V+;��)��bN2�V[��ɠ7�u~٣N0�?b~�z��U=3j� ��vr[p�;�I�K'��n��4�l_�u:�tP�Z�	�!��L��b%^W��u�)�c���,t��%�M��sW��e���F\����d�_�}���&FÎy�]K}�����ܛ�y���꧑�Z@X��~�l�%~X�B������v�	6�ꗾ�Z����gV��R�풣�����wɯc7y��,t�Cxa�Eb�ncPː��W�*�\Է$���_�����H�6iŝ=	��P�.���MM3�:���3�V�qh={���h���x� ؈����_Q��4�}�V���#��R�2s����)*,d���&0x9k�x��f���tUR��8=�B�U���R�uN��ޫ��E筈Ŋ�F�_dP|�x5�֣�F�s�^Ξ�~���U�1�Pē�M-���[&�C���mk���QX{yd��C^�� f�`y>a(~��r���>��R�o�Q]H!�^�iP)*W�C�e*�x�~0�*T@�\A���Û��%t���f@(�!(w&�k���-Z���@����5˳��kR����i����տշm`:���n̂��#$�W�w�{�v��7�"�
d���Z������J��gӶ�_�=f5����%����W����7�e��/7!�0%�f�K��Y��w`u�	Z�`=q��_Vx�W�&�[�
����<�ǘ� �]�Nd��/�S�.���[��x�I���P����Vg4�R:�v�CU䖙�*;I�**m�'�nf|ǯ�������cg��Ssk�y�Z"m�i��������_�s7���&jɚ�W��E.�8��A��4ƁN��.�~|�j�*�����N�u�Quwȧ�ȅ����S�rZ݁+�3'�oY���d}����e���wQ����	���8ܧ���?�b�Q��j�>7��ڳ��;&A��L:�"3��N
�2�KF�>�9��E�JA��pz0:�Cʌ/�ZZ�3��>�w�JP��7�W�'e��ߞ�B��օ�l�&���y��$�E6gƛ�7j�D>/�����O�����,k�my^��*Fw�1mu����u�2�U�U��͡�ČkWp2�8M���d��W���O����@��+1�7Ua�Q����;���I�P������r�_��\�u�� !A��fh{Yw�9htP�m)�j������rY��s!��)���d��0���<.�N��}���bf��@����[�x{�#XG%CiN������˔lª�H�]�INs�\�ꅽ���y{�GM����X������uàb �5i6���z6G�	-|���G��G�y�݂�2Q0�pN��N WR�
�^�n�����w
����r�^�;���eL�qk��岒n�'������p~w	Ƭ~� �h�;T���/|�����ܹ�c��-�+o��ޔB��IZ�x�4b�X����a��M�*��PUv�+P���}Rƻ�:HU,�JŁ�@���p<������,�����ƛb�\m�L�~Ҳ��h-���tH��E��"ld�4LjL��p�8i�����:�VN���9��uB9�3 �a�%Ts�Kq-e-rA�����O�� P�)CJ��r�lHOy>n��p�P�0����dE����t�奪'Y�|�PJa� ��I����T�����,���|!�$ l�B��r�Ϟ�s���g�wC9^ו{/'g��E<�K���I39+{����(\�<r�� 3�JR�jS�h_+��g� !�|�gѾ�1�ŜF�r�j��\�1AS�'!����[��(`��#�.KD��ˠ?�	on��H�B�n���v� ��5d��c�ऀ���t_��eW��k%SqH�S��Ypv�{ �t�F)�h�֨II��<82�:�W����q�l,	�s=lo���5�Z�e~��zf/�"6��(�#@����uz�~�����]+�)�{1��7�s�!�5��D�Y��a��PRp�o�s8=�,�S��`�wkF�����L��m}��: I�����e_{\��"c+Ҡ�F���!G�W���[��˩����ͼ:;Ϋx�����{�l
����^j8��p���"K4A���9�����Qp8�mE�X-y�F奂f�=���n�d�������	u�>�	_`)��p��fl�hѩo�+�%T��C�,����|B��i$LD�J+ �N���=i�F��⩔��<�U�S���	3ڐ�!]��d����Æ����b"L<C1/M�������ɦ��C�o��<K�� *��6��LX��`�\��̟i�-ROG�`&�u��;U��犈����͗L�k������(��"$;��$��o��j|�p�gB庹f�檁@/�;���d`�ln��o6��@�Z��jܥ[�(�	�o�#���TtAt�s���v/3�Q�3I�����g���dgi�z!����|�c�
�;֯M�X���B���~q��>�����w-S���������;3����M��޿�PK   ۍ�X#�@�9� �( /   images/bb1d7dd6-69b0-4e8d-a72d-bbaa9fc3070c.png�eT�m�7:��� %��1��t�twH��t�" �t
H���"u"%�Cw
C���<���{��q�^�B/�9��<�w�y��&����� ��ܘ�@��o�;��R�pݥu���?����-Cw����a��nއ������^�nV///.['{ws+.g7��m�-DQ橎w��O�#��{y��	^�����}.ߡM� �ħO���g�M5�ޢ������`ʝO������S)C&�J�Y�D�MCc�6݃�䞿p��i��A����m_:E}�Z,Ho�F��B!�g�!�W��ʐP%��y}�3�G���k��v��I4���f��뿷ŤP���ƃMa��z"��%ԙ.x��l��?����_��,���9���mN?�,�#g�ߚ�D��ʀj���� wm��ߡ�?L��s�{�+ބ���}o�-�L�4'�;mY��iD��o�q ��Z:o�)y��G6&�i-P��~B뜰(��/m�a#���h�h��!�:�6'�~��Ja[�.��0�ū��|���1������.��=��� �r[ f;�VW�GI���r(���1'e�G�
�6a�@wq��)�{�uc��Z5ʿ�k�g���$�Dx�{�e{�H寞�8��J����3m�U�P8m>&+�{b�~��"h��T<�s@ �X��q8�Ѕ=�XxxW.�⤊Ʉ���S�}�Љ�4ߊ��R�7�1}l�y�ͣ��5g�U�,� �'M39j�X�+�T*t� -�#���KB5F���\9�Ϳ�=��q��6��:(.���<	�&����/~���
ўF�\b������L��NTvw�%�h-
`lE͜�"R�� ���	�zS�����u�rL�����v�ʟ��r�1������	�����_�OKZ��-����D���om9rX��Ĳ=v��K�434TQ� �'����(Qa�J��ܵ������_{)W��V���=Lxҁҭq��0���5a$+��]�0pȵ28�쳮���t8��cbb2;5�mt�\y¡�f(K֙�(�D�y�6E�A�i���q%����^^��}�&��/}�G6���T�	ŝZ��G�*G�9���F��Cvy������u�Ү�<Ĩ�!;�Q$}��^^;�����>e�ͥ�\^^4�۷�v�1x���B ��O�l��t��d�F��=�ä ���l`5F�*5� �?X�!��G��r�.�
0̜s�*�Coa�q�mA �4��{6�`�)h_�K���a�C�l(!��m�|95й�{@���y�}��a[�$�UsA�hc{��y>!W�FM�=v%1�?�F����$w�c�c:�H�mxr2��?�k����\�y{�!3R��V('Ä�bC��C������A 	[��~�M��܏�����p��:T�
��c�k�ba���1D�1���ȝ������װ.�x�8�2��c _����y͸����\"�M�z�G]�\�|Pp����m)��z@ޘ��⿨����Ç-OF�'k�Kkkk�?	<���<Ǝ7����7](��q-�b;��~c ��
�dg���K�;��$P�=�r��b.l�� �=�9�s��:��ׅ�����m_G�m�A��.6�ׁ�+��|q�ݦ/���W���P��n����m�ԝW�t1�&�Q���I�4��s��3i��0n$�:�L 큟�a��O�m�>��Oؗ�WnBn�מ������G��ֹV�54h�0�V���2�cAZY�%���i�3m �����o��P�v,�sHUv{�Q ���04�c�p�l�8.�(������
�*��H�}m��{B���$0����b�.!��	Ʊ`�4���+f�ؐ�-�y�4�K#�&��A聬��Y>����xY�W�3����aH�Ѕ4n}XI��I�p/^�e�Rt�tD��pE�U�6��9_GW}���/��IX��K��������/��=ML�o�B 5սk[���2�T���Vg1�ߖe=عR���j�Ɣ�����hxU����ӞtAw���RxE���(�3ߥ�6$_'��*^�o�gN+� �	������I��'$c(����k�I�o�I}�6�]��n�Rc����U�r�"���o���ђ��ēY��J��ã����1�����P�d����2߁��N"����<�(��Z)E�;>Ѷ;�A�+_�w8��*�g5v�T�
]_]�M�Rq�ĪK��IIMe��"Z�_I^-
����hR�hY������(U���J{��DT^=X�;b�� L���Ԃ�Į�{����Z���J�k�+ÙҘ�����r���2��0Jj'gf��<�i8Z]YhOa�����y�(�"��%/}��w*�R���+�x���~�t�-�S���AX�J�>m-	��^���_�L�S%�C�hM���� ��.�8����۵��S��/�gGп��}М�ѐ�k�cR�6E��y
Y�e1Y(5gQ�B�>��[�B�H�!*@�}��w �d�<*e/Ψ�.��u��'8���j���U�Ƃ�>*X͙D���U}�s�Ѵ3N݌�ۇ�{W#��^�${���׉�}���Y�(W�£��?�w�d²���Eg_�tW>�m�=�J��nl�A�����]�g���
/ߧ]PX���/��������V��Ҡ���5k��T:�]j�xl���+4=�g�~;Ql���h����x̊��9j��������q��U��=�_x�����_<�D9E�ce�v����㵤Z��P��&E�U���*�i'y��;��1���o�u��y��zx�����s�{,	!�Q1b6�@6�9�1E�0�r����.��)��XNBu������>{�_T���Ao�D��u�	����a� �Y��1>�w. 2�X}˚��И�^�BWĶ�K������bt@����fT��s���2i+����G���$������8�6LMj�;��{
w���s��H�X0)j�\��䰒�tX3�2�g�FV<�4�S�D�~�\�)H�׌�����8����M /�7A����&�)1Y�������)� GcÏ�`�hG/�-��TV\|3U��ް���2{�������g/s�L:���q����h1������gK���OV4�s�A8���؆H�R=��c����h�8I����J�vmrӽ��)29,W5O��)�]���8����O\#�>��"��O8�)'p�-�$$ԑ�c92>�g�a-B�["ٴ�N���,��3-b���DiQlw�0���Zá�"�m3]���閟	�ۯ�c�3O��>B�nܶ��8�w�+�49�P�F�� ��-����x`����B��'��(N��.�?���rj���x 9)����Θ-Y�L��s�:��Qt��KH��Y�{h�i\��XHBh�y~�<9=o)ݪ��?��Bd���\��	��F��-��Ԧ�~ͣרCs\���MV�od�u���^���G��gQ�nR�A�Z��tĐ�L<J"X/~rrp+Ξ��Sl�gQ倠 �i�,���+&b��a�x�V�`�x���R��6>Tw�_L���\�Ɵ�y1k]�=5��Z�L�	�q�W�����Ó��ʉv��D��<~ܷ�a� n���ԼI�FU���T����/z�K����G�1�>��+|�S_v�&YGF6{��t��W��/��*3a�z�z����򰜪��3��4�z����N��Ϡ	b"m�2�Y�E��~���E]���=��g�+R;�X��+��􄤯[1�z��|��[���r��+{��Ɲ��ʀ��\y]4A�+A��φ]!q�4��x&ި�f��qW�*�1��.�'O^��p�+qJ+5��Gu�Z��Lz��8�%^�C7��[%��#��ޝs���,��¹ C�˩Rb�逢?e-*��s����>�����4��s+�6���|�����]�aտ9Q�o����`՗�V��5\5(aO��7ܰ�`7�1�'�ӄNU�g5��~�7p"��oBk3�kNӱ���9<��3+�r"e�޸N?ç�rE�Εs �xّ}s��ƺy�=���G}���8LĊ����;8bj7t�뎋{�/,-�Ə��|^?�C��ǻ��<��T,Xt�O��K���怤��t�w��"�Y,Z��C �M|��}��WT�Y��H�k�%rBs75jHT=�9�M��%����rnF
P���}XF�
�y_���3yV���j�و �.t�E!Tn1�[{r����hh��C[3�وA_��AWE��Z����YW�	�R���?/)���H��g�5�{a#ڧ"^��g}���hO��E��D�U��_ʔ�r�]Xs�����_s~6͒��S˫�k����z����z���-�\� L��ϟ91���"*q���N����EediSs����H酡j	���G�e�%S��,}�KW������,9.��Zn&�}	0� D%�2��W�����$l�$:��0uj����j�[;��z=��UKC�gX��z6��L�Z�F�;�c��{UѬ�ߝ�}�k+�RN�n����.�.�iy�%�,��Q9MSX��G��~4���7l7l�����p(�zb�N�j[JF��c�:�){���zr�6&�� 6�HFN����L�����[Z�ȸ��꩜ͳ�nՃM��[�HV1�Bz�Zm��#�+>��C��yO�˼�Ae��8��7����Hao�.X$;��e�[��5�Gk!�V+���gA���9�	d�4٥��i/�IǊ�f�S�:*uT̉}���q[������m�Q�������� 2c 	>5���7�s]����#����Zn
JV��"h�gvPN�
�"򺿗�k���
K5A}@9��u�f�װY�=vw�`�wvQm$pc�PY��a_���oYf���V�&��%�PJ������Lu6~��o3T�Ǡԥ���r�v�]L��l���j�`V6��$7��?�8�+ye��=<�
�J��x�h�~Y��$�B�Ln/b�E��Тs]���<�5\��ʶb�:�*��Cέ������W� �f�hGa2�� �=�|�T���x�S��P��َ\
�MtY`z�^�&^�D�����d/� ����!s�	ߋ�q�.�W����Xm�l��E��f�Xo<{5ܶ<�6�R�(�5��?��Gc���-p��_C�^Z�?j#����Tb�ڍ��Dd���7޾��V'���~��'���pj�9� ���s���:B��\�=�HS�Q��76zF�M���WÚ�6�L}��Q���Z�����nAi� ��07w+�^AalK�w�.���5��T�8�B�����g?����:����X|��ؗx��N�N�/-j^��COf5.��A��i�疼��3$g��]�ѫ[��O�8����(�Hg�ݣl�0��,�����"z瑞G�]�g�����nƉ�Y��C �񨍿l��4C�ը�	6�+���0ѷT�5���2�xp=��*os���u���o����X���>�1ab?q����5d�W��������9�&�v�N^J��1��.�*�*��I]܈3J�l�;��=�1� �}�F�Pxv�C�U�x�:ߠw�XV�?��y=ξ�m���&�i|�P�]����ڨ������ۼ��sl�]�'��x/F�}5D?�æ���ҪO�&L��ڵ��L>#�4J��a�'��"Ѯ�%���s���߄�-�g���x�_��.��o�a9#�T;K�K�!:�S�?<L8M��68<?���������/��]�ێ��UƩ����Xp;�����C�ި�{�t�&����8�y�H�E�Ba�Qea�K����i��g�gQY�����ִ���P��B����<A��;����\� ػpcP�
�c� ���aPMe��C�Rf���}Tl L��,A>]w��E��VX�^`��H"=�T:LJ��0k�aP,�/ б��|h��:+�\P��z4�|�,0���f%��	P�%"�٫w/w,D�5x�;q!�w�Cϐյ�|�����>2���짿����֎É�ප4��n�5O��⥫\~)�!z#U݅��GI]��D�����cT�-�NO�m�c�SXR��^��JMM���Y�����C,�ky$����g4Y�$%"�P�U��'���\�Y2��,�����p"ڟ��)�!�T);�~)?���k*⢣{ݠ���,�a�s�Gz��|�^��>���)2����:��ց�����������Tg��f;�7;pO��K��vh���EUJ�1;��H�b��~Cǯ��/�^�&�w}J�s�+mh��$d�';L,u�%yihՕ��<�	�T��<M��Sd0�¨K_`m�9��~}�ϛLD>�vu}�ږhxb8��PR��5�\�4��C 3��vk"�q��W&�h��O��ԕ�w�_RF,�0�J������W�k��h�S�S�s'�����^+�MX�����ǵF�Ln��lܴ!и3��ܣo�5njjR1�����1�jo�q]L�pO�㝨��&�Ԯn���JK���8�Z���_k]FE�(��>ܾ��$��ח�ä�%�������BTMU��0A��YI���Ok"]�����$�/7�@|��<P,���"�T�g�eeP/Qu�l�*�JW+-�<4�Gcm楓V�錫x��=�v����4�x%�[BJ��ӊ)ɣ�R �ݔr����"�������Q�j�#
��3j�+g�{����i�V��"p�¸	�V="M_'p9U�z�Z��j����@�B�Y�\v22h���Ͽmak���6!>?��ޒ:�تȰk9q�����EQ�k:�h�[Ђ$���S��;�%ϼ��4z��4L0}(< '���oC�<#z�,W���Wx��Y�;� ��.A�v����<�'=�!~~_$����L�9�~�����Ff�`Sg6��"�a�a2�p\�O/+�����	�2�{����'�=��/�6?��5�TH���z3�E?��uUf$�Z �H;��b�ƭ>�Z0��Q�
�䆅r�e����&Ƚ�.��'e������,����mA��SD�fj��XO��d|�������O0����޳��j�����r��O8)l��z 2�_�B_��Sl��=�LU�2�IS�v��qhy��,bld�lѨ��lrP??��������cj����.{fr�v�b~�K�d���d�wƫ0��C�rs;�f�B!��;-%�~�����㿫=·��nZ_^����jEJ��e�TV�
B���Rl+�1�L�G_�틠$.��yz{�^E+����0s��o��x�����2�1�:+�Tݕ�Z�}+=Ƭg5��E�8Z
�q���ҳ���,l�.�kB�-'�ř͞����_��I!�/6Q3-��Ӳ_;����fVIz�V;����Q���o9�z�5�y(�6�\x���|W`ƣE�A>�}��L�.UPI�:����UR`.B"�d:c��F��
2��*���}��(�V�(��f��+J:~_B@�*��&V�bj{�6#�yV��P $��0"ۘ�FDΰ���=�h��琛[���Zb��0
^h6����9�Ų��i㕠��P�R���g���I(i�0�V�� ��6�>j+�h�~�!�����d����|�e�pK�Rv���q�H�%��<��<��\Z�~�v/X� ��"S�1��x��!AKX !�Q�{A�QXR" ������I����c�vv�>�"+C��Y!�j��5��g��\:��AZ���k։�LsI�Lg|�.?[ba^���۽�)SM}��o�Xd����Ìjr�"z���b�@�y������; c#!RQ1�WPl��zme@���l�Λ��������;ޡP�{A�>�H�Z�� L��>;�ä�Bw��
�^4���l�?��|�Ǵ!��1GE�Y+�g����x�d��I42>���1�C��Ç����hI[�S��J/DH�V\�"k)��.m)��as"�oG�����@q4K�[���m�)[��X���)	Bt�̜E� /��s\ʄrO������d���S�=V���j�qF�X:趉�~����]�~���]�A�ڱɃI�=���P�1� /�oڛ�&n����
�)�W�qK�GY$o1U�W�4K0UZ%4�|S(��uєif�%#4+&���#@��<�͙9�����C�n������x�'��n(eTs酂�|,J��:�����&��Y�yr'��
��w1 ��L�@@��[�}$���D����V�q4B�� ^C�F'��K��q^�ܫ����[��u��e�\�V�<f���},C-%�����ū�W:��3�S����g�>��Z�4o����?e��f���K�[n*8X�X�/� :H�r`4W�+�P�{^�o��(/{WXฎ�{IB�i_,R�?6�����Ǐ�8�+p7�@=�R�&v;��J�>��~�� ��G��}>� �*]���N�%�#�a���Ɇ�v�7�)����HP|�"vx~^�����X���H�Q���^t��IIb-��}>?�l���C5M�`��qէ��&�{�*�ؔY55z�S.ouUyV�0z��Wq".1W{���{>ʏ΄u�y�^Geh����\W��ɋyi+�m�+�Ǩ�EC!�YUs>��!����!a���
i�3w�������I����ji����X'_�	�<�d�D���#׹��D�Lz�����IA��7C�s�-9\�L�^��fi�����UR;�q��F���	<��zb�I	���w���O��0���%ϰ���v�=c�^O��=�υ�j��V|@�/��Q��F���+�uA:_�c�g���R tr4`9=�,E����]�����ь�3�)^,vG��X�gV���+貔��K��ʏ�[$k����~*��<;S*^�k���?@s�"HI������V��7 *$gQ��8L�s��ĵ���l��<���?䦽"�ؗ5���u{����H����jE�s�Y�������*�s��Zl�;��RD{������1�ֱ���'�/Y�	�<?^�#yS;m ,��mOn���XlWC�z|)Ѭ�}@X���STX�+�U���}^�Е��{�"bB�݇؜Q��`�|=��Eە$M6�lO�ݖi��3�Xh��Ɔ�Ǻ���� ��fE�v�qM:Ŀ��#`];����|���U	��+��T��  �J� ���m���KB(�?�׹Z� �G]�\�p�����g$����3a�/��̃!g���Bv�׌O�|8;���;:�,�c[����j"=��� I��J��6»��|��7Vho)�����
�[�Ұ�Ӎ�O
��o)��׵�:��wAtE�a�&b� ���kD��e�fR�����Ll6 =���k}��DzC�,=�g������ ���}�#SSŎ5��̃�;g��"D�~��ғ������>)YNsfk���Ѡ�h"�bI,��{�Z�*��q�vT9~�H$3�a������Ҳ7�Ud�#��i�IP��fe�o�R��J]x�ݨNx�eM�FAQ�0h��7��k���W�"��=ۙͨ�kOM��n���j�K/���GZd���f+bc�͛�S�&@{��-�	��`fr@��]ZXȦ�¯8==��g��鈊U`��uR��N{�=�O~☂TME�������S��U�0�`�T`�k+�d8��������V��{�Շ�-�5X4�A�o���Vn

�q�FM�S+���yPd��@Juz,����o�	��X�TB[�=�1�9J,*d��(�-@����(�0o�d���EsN7��_-�r��BšGE>��$��l|������e;4�z�2�y�W�����TE$Y�xP�W��H��]ݲ��KgF�]����ۊ�rي�0���6��A|���1G������{hJ�[�`���vo�>xE��'L�g�K04��v9��l�����e�G���ŕA�5���g����5ԽT�ۻ)�DIi�Db���f�)�`�{��O�Np���R$���^��N�dR=ƥ �b�k(���M�W3z���EԊ#Ŝ�&�rN�V���3�ws�%  �#*zr4w�lgOhT�>\�ē�s/���ɢ�^P��G ikLQ�}��d.�i ��< ��*��n4�����W:��t�x��m%��.儭 � w ��bs]��+࠴��ݯ�ǂ@�BD˿�vkޠa��#���[S��뮔�BO�F_G����$�?k��0�5!&��5ࣩw�v����g��ڡ�?�ή�=�Ѕz�?p�Jκ�B-�9ˑ��N4f/j@�����dh���m�Z㢾�F�='[���U�͓�����)��//5�7�韋ҩ�zӺ|#g������G�Y
b���,�b{��^�U���p������L���H�.�1�ȅ[��p����XE�Ο�f-uqk���9����}�I�<%xgM�svK�(�hgB�]6����v6�db?>����9m��Jcl��< {.g�TQ3���"7oF�x�k+̸��v�{�	-kȗ��B��g�?-A	�M���
�y�_�w�#@e��l�OO��h�h8r~=D��x�\� fclD��(k�t�xyw���s�S�*�
d}r�:r`�{ *�846�J��R7*cF+_�,�7�N1ٮ��Q,��y�9;a'���L�@BDw]�t�q_���5��EI4T��!����B
��V
��s=�69j+�����a���a3��G2��C���ё�_p"���Xыv�Pm�4���J]C3���Q��>g�~�e���s���ܰ��Q�U�������bB��{&(.��˃�WX�K�)ۣ9'4 9B�-0�|�ǳ� �|t���J�A4�������3���٥��:��f&b�����){�+���l�*��Ymc���C�t���b��>CZ}y�?�/I?�C� ��&��� p>	�kO�=�i�b��4Q5R&�;���+3�Dks�J�ti�n�F��#yT������3`^�牛��֨)9�=���:M'/b�3��f=i��󰷺:V���s��L����Y�Ă��2U*�� 3&r�A�	��R��/(�m8�l���!��{�g�3n����v��n���Y
�=���K��@8�?��a�ֺ��[��χ͖F�������Ο�y�<UK�>@N���u�,��\���5�D�ϸ��P��;z9�-6x�3-�ė��}&�dӫ�!d����,a�ޠ	�����]�{��z�Y�M�`��y�����dn�ž�љ��#�_f������r%Mk����DʙzgZ�Ps�Q�t�J���[c��Z���m+���Gs�׳���ʃ��a���"rK��J�~W�\V��$�91gϴH`~��
�Y['��NN�n����vqr���
m���8���c���=�a�F��?\��W���x�!��ST�<���p�?^OKF�y�x��\�YG��B	<��q��^|ZI���i�U,��L��Eq�;��;��{�#�d_��!Ò�s� nɲ�@�b���QmV��l*f"G����"(��Fb������6�~EϹ�R� �L�O��h��S\�Z\����gk����=��@�ʊ�z�E��[�\�A��+:��������$��W5
=�����M����Ua3F���k���Q�A����c̆o�1`��MԮ]+f@��U?��!Cͧ�G��|y:�ją~dt��i��b�iޚw�nMI`��۬��&h��1��s/�	���t���,G=����\4{N4�e#%�C(�t/���g��f�
��1
h�$���j�6̃��O5��7�4��LSR�Z��a]v^^ELT��<�k(4�X9��kZ,��_�[���_b2$l:^f/�=��IIyr�\Z�c��*��V귭��v�/֪`�/C�kK�����q���M;��An��h����sf�$e�նI��W��Dx��?��f�K*]R<��A���޹k�Vm����YU��}B&�ڕ!<��L��9�O�S�}����X��ʣX<�J�T*T2�`��/W$G�S�[Φ;���3U�J2���B�k��k������T_OX�rMU%���% n*9��Bg����3�M�p�HF��)�6)��^���>�,٠�;���2���U����� ��JN�{�"rs��U?���Rg��g�n�\O�Eث��7֟n91f��[bX"`&�c0���^۰}�\q�:s������-+]��e�"r�9��&%T����v�o�
a�+�G���j5[�;e�A_�æݡ��e�zۜ��������S�%*�����<�(�Q�4���i?c|)Bp󧉉��4���~�N�-��y �0����S���;�[��<�sr*	����3��k�F�X͕������*�X��T>_��j�;����fN!�a���GfPR��^^��^�~\��{�kRr�+�J��,�t�ǰyNԊ��=37L�估� W�dpY̋�]���ł�Z��;�cV߷��ci�nE�)��
c����x�>%A�$c�S��b"n�j ���M'����������j�����u��"�J��u�@��C�����b�z�s_��W��#���vu(�f�'�e&�\B�[�ɘ�������{V�������LC�d_�C����5X<�YM�lD:��v�8sFb[���B��Q��xr����T_�s&���n�S^ޯ6�-��4���&�=#K9���$O��%�;��v]Į����ɟ��g�s��Ν�GJ"�}�3���{ɀ�yW��屿8�l�?-�)T�L���܉ wn&5����7�]kd�P�}����r4�I5�<��?瓶�<�{���M�5�C7�3!�E��+��R�aE�����%�Q�%�\�1x
H4��w�쁭_�ڭx�u��J�?T���*����꛼�U������%�5j҂�&�L���L ��)X�;|�
:a��*y�Q����p;���_�a��7���(�ϸ�י�d<C
��<���qGT�J3���`��#�æ�7k���o\o�]�oշHs�&#^�D�O/=M�|���U�*m'gƌ�����w#H�5��^��gʾ��6�ʋ�^�>5���z�v\����Y��@G�Y	I\��N0K��`�����T�I��������z���f����@u��ޑ��"](�{)��[����٫_�Ah����Ŵ�2�$A6m�2F�R��ܭ#L&���usWo�O=cFT�kUߩ���^�A��9�*�������z9�U��!��(���7/9���|NU�1������><�(�S�:N��RgW�i�����Y÷���)�aI�����@c���ـ���syx�	���Rm��D�d��/@);�z�U�pv�$8j�/_���[\�11#�x�A�axga��l�z�1ccE�H�h0�����K�=b�f��@ݘ���MJ�GV����% "&���,/fZĪ=/�g�����Kt�O1�]��9��U1$�r�m8�F2@�_������\���ۇbǄ��)�c��?��x ����-Uc��I٤G�X`�H���ckt��o/�Q/,����^]��L�w,NK�Z9�\1� �;�Ub\�?���]�/�Xyj
�8���8-u	d)����~V�&�wG�#�D�<]�G�öt�i�۵I����mj���<y)����'ܮ9��^��o�	�����ʖ�򟯢H�Z��)c��G�Rrե-j�W����9e��s�K�P?@L�G�X��E35��C�]��+X�%:�����8�����L尩X�u��i���ˠ��m�e����^�����k;ӿ�3�I��&����5��=Ch�V��6;��6o�6Y@^�nT��6���-��[z��]����-�']���*y��I6b��1�e+HV�ԭ��&:|iBDσ����z+G�`��	�������M#�׉e�'J_���#5��ܬ��?U�j>��k�#�Z����ʍ���re+ѹO1%K,=�����+����N�]�ȷ�[نު�xo2��]?mB͂u��t���.�»L�0-7��N�dJ��"F�0�B��&k���fIB�縲����Dw�Ȥ�/jq��y8�%�\��a�Lm�o�x����-��(�nn�K\Z�����Ȝ�	�v�G݉9�PC�<Q�aⰢ�@t5+=MzP�,N7�M����r�pP6W�"��X���_L�r�k�Z�!׆���H{))W��3y��LF&NҠ�<�.�4�^�|�בm�3��*O��hF���B��a"��'���(F��mW��w�~3U��,#�ǛXxk5w����ǁ"��]Z�"������KQ��W��A!�!���^���^����(N���}g�f��U~K)$l����A�w�m����s���ڕG�{���Ʉv����{�Bj�ƻ;�>����a�+x�5��<��o�?�v�@��l_��ƁJ����P#��CI`sl�[zft��ď��e�$��<w����__u��D����f�	�R���&cI'Z��Y�ZV����ż��~\s�x�߹}>E�Cjw#:e�i��8�Qj2�?E�K�n��᭜k��ϊ������O��7R�wo�_'e�Ժ���}:��5,@ޔZ��i�a��,�~Tg�FJ��b��&�hޭx�qE��k-�%�]h�G�RT��y��B|�!�o,��p�B�k�M Z��@s����_k#u7#0>)�^r��
n�{T���R(�K��;������EY�9:��殆���S�*{m���X~k����b ����f�����*����KJJ�L����x˭�J�'8`�ߛ�A:u��.�����s8��J��~Z�s34f�K���eJ��RY����ӎ�sGy	PˣU%��enG���6���c~z�b�J���g;%��&�φJ��<����V��P��y)�f��?�x���s�	-h����JW�מo�E���'����ѿv	A�媌OQ�;�����jI�1-����p�+�f��-�^vYy:,�:e�#ŻP�.����A�)��^���Tc�w���]X��y%�n��ܘX�\^�i�|޷RP�P��n��`�;��:�u`��w�.�@�D��`������v��Qa)ysU&s:-�O��E�Q�j����	Ґ�>�9�@��0B;����*��Y�x�,'�y���n~P��Kͱ˷/Jު���H��^�=�(�g��4��<M14��;H���@�h�R�~�J�b�_��"�zn����+�8�D���M�}��O���m*�@"(����Q�;kJGT���C�4���4�&!]�	=����-5^�q���5t����jF��a-i4U���	˗�o���cКLc�L}7�ŋ+�w��p�^�'�!N/zӰ����D�TQ���!���;����t�(L���ň�%�n^E���ն��vb|R&�6٥a(�E����y8vn��k�*c�j%ѕn˻�,�גWG|ٯ��U��Cq4xZ��BC��a?YE�mi��~��p��]�kep􁿢A��1u�r��<{_���Ú�<�73�=c���l����-���qE	wN�N�sh�8��Z+�(�Q�}�*>�^�̣���{22���a[Y��kQ�,.f���A�"��:*����le�<���V�d(�׵�sZ�z��1�l��9�rb(��m���c��v�@0��A������옍�<v"R7���zbX�3Ğ�)~}X#@��0�jV���hz��l�k��`6s����@<�!�nZ��N/	�������\j�t�z�F��n̄H޻e*;y��r�*��Fjq^k��C�%Y��e3 ��*NV��;��i�em�j�W��vHV��a�i��i���� �!�h�-թ���?(���w)m�7 =���CBӨ��	C(����W˒�Q����}E.Ve a�Z�����*��Uai`"�I"�$@k2]��V�e�L@���'�R	"���4	�:����]\~�Xm#�h'�GD{Y21���*6c+x��v��L�80�UQp!�"���ǹbg-�1xB���L]H���-a�P�䙪;sI��cƍ!��0KA�-2�:n)��ʵPa��ؼ����w�]�o�8�p0���)��;t�GH�7q��+qQm��Y=���|���K���hC�������a�����л�ب��7�3�p�HĈ�e�Waq�-�nW�;�hu�k�<��1����0,�������=�ݧ���4ڶ�I�ʓd�����F�&�g�� A�]K
��w<�ͶX�08%�݉N�ʻ ald(���$3�cRݺ���"�z?#z�4#c��[%|ޯ�F���Ƌ�<����S|�M�J	S�r�6�	�Z�/Jt�E�o����47�� X��M��sX󁹐��	�B#����I眀�g�X]$��5dRb��Zn�t$}�N���C�Ljs�tr�Z�����w�:p"���Y�3X�>T 6���f���ROȗ��]�H���vU�nK�w�M����qBZ�?|�NÔe3oЗ�
��x`Tݼ璗7�%O�iхr96F��N���s��q���OJ�u�s8����ޮ�9[����r%��>�߽֞{��;�qRT"e�:��L��[�P�I`���d�"�����,���-{!��p��TYR��Z���2'a��0`��ӹL��te>��}3|��^� �4k�y84#�BI�Ϛ�&����X7L�̐��9�5;���>6�1뎢J�] ��5����T�� _�q��.�v���Bߺ}�'����Ng�\%o�u����X T|�����,����S��3BW_1��.վ������Hf�����F��.�8�(����R�k/��8��_BEȘH$no���ʾ�6����ʰ���m@���G�;�C)�)AJ�;��!�C��v�n$�k�;���^���8^r��묽��^�Ƿ{�3��Z_��ûhˋx[P���;�
I�Fa[4�/ۃ:�`��n�84F�B�ڵ��x�����V!rž���Ke' ��Z)���%"z���k�֑��u�������͇G&F�^�Zi��+�A�_���焜F�)�(�]�v~��Y����哊`b|Y�������vW�>���T� �)�O���W{��Ŋ�ε;����GeWヂO6���h��?��O_g�&$����*�c����w��K�Ƙ�<�8'�>e'��Ԫ1̦-��2ٱ�%v���g�)<|%#Fr�ۥ$V�#���[��~ڑaJo��>�g�Ye�٦�q�W�d	�~�|���|S�č+7 K`�n7�
C݄��O}^J����A|{[ڛ�ޯ�H�*��;r�b���fGU�<��2�y�C����o�f�a[.��ݣ�Zc�}N����`:�jsLv�jE���褷��3J��:��wM���L��D�p�]�9��ͪ��q�^�����Чmb�#�T6
��2"���&�R�� ����U���rD���e�-��Mol����oG�Fj�|'{�ߢ@�7p��Ch*C��h�r5��f�K1�O)r�L!Č��K��		�L�2��8�ؼ>G+��L�+�F����x�����O`D� ��D�6�-JR�h��=+T}��#NL��/��|Ig��Q�"�XH��GsdL���
9+C �X�i�R���,�mx�K2�NP�k"R�`���r�·����j��g;������
�RRRmw���DW�D!��RU�-������t���W7R�X������,�����l��7o��ĂU��u����\ O/+��n��
iR���ڝ����r��8��h���g����`:�쥏�̠6���"]�X�ו�(C���?�;\���8z/�f�X������ub���i�k ���~���l�����8��p�h$�RTûI��?����o~������������]m�@ۗ������I�\�a�\�\_�%W���NWi^w���3V�̟K��ׁy�*��M���#!��u�u"����;ۄ�:�����B�S��S���W��g����H��E�Ҿ��d�pb(����MMQ�Y���k��V�ƿ�ao�do_ޡ�q���ޣ��k;���s2X���h�k%�|�C����J&a�x�P��>�f�x�p*�����Zk���4,N�&�k�pg\�,��V�Щ)�?:�f�x����tc5USV;��t~	�~�S*�X
�j�ڦ������ęIi��	���/��]+Nt�0t�P��r��+s8}rW��G�6^Y᚝��2��[C��O<0�Nh��2D���:�;���9ܸD���*3
%�KU�[WW\��)gn+(�)?ᇔ_U�(�2�J=�K��Q$n$��3}q��G�F���{'���K�����T���~,[`��C8������fdTT��������
/�U�$�	R�=Ec$z��T�b�mն�Q�&�̮&uc���t���� 2%7� �����W���脏įY SL!����������t!JQc�~��E����"��<@5�$U(��w��ڇ[{O�����!�و
c&����=`5��K|�� `O<zxl�p��GK�w�_c��-�C�4?\8�����S[����h�� �C��)K��k>0{I��|'�!�;����@�\8��@� '�?R�#�d�n�
���/*0!~��[��ÃcȈQ������iX��DG�:`b���������� IG
����0�~�h9�������?�ATJP��o�HF� $����J�����g�W�j�'D��� ]��o�+݃�e�#�*��\t�L�* h�����GE9kq�߿����������'��B,���?���o՘�k�|X2���%K�FT�.�������R��Br3�QG��Z��X�k>DvB,&��.��Q/����j�A,CS���q�Axp��7�1���aFħ6�ߍ�J[���7��Ӷ��w{���f��u�+U	��G�T��������� �n	�h���m$_-�&1�Ě�1>͚��cd�2�j�k��uY�'I��{5�w�=$Ց��,)(��

�U7J�\- �02��#$9E�:�vW�O�!���d�A`�h�:�Z���ħy�R���^�k{� ��޾��2�e?|� ��ٹ<�gaHк(�D�ց��"/���b8�0 P-�����aw�ſ:::N��:N,��ߴ�X���<�!_���`Uw���k�`sB���k������[l6X�Λ�	>X�7�%%���/�W˜י <f����P��|x��U� C�БckH:������6wM~K�� })Z����Q^�M����M^��h��We��&�T/n��G%�"i�Qe�)nsrtտxj@v)�vq�7>�&m�*��jCL��������}{���}����:�ɪ!6u%����x����CwZ�ic�W_�|_����h�%����Y·��(����>�{�4|.vp+8>'cd�r{���Y����u'Q���[u�>�ܓZ2S����2�Q�. H~�˂H��r�>>��ap?���pLD��+��������՞"���0��Yh����+?1	_Tڀ�hSZ?嗹~L&XM��)���\�������)��Os4f�q�mB�O�G'�����+&!?��/�iٷ� ���<���H��:0��>~��_e����Hk��񊧌�e���(�V2~=gUR��N�V-���e]�~̹��W�+��M7L��:f�b1ʣ'��ГD��W����:���/���JS�)�/��
�H�I�/�y,��b������>���;���V���0\��؝Ќ�T��}��L#?�.@L����Y��� o�LPz�idP��zX���ib�a����'Ϸ��MYoE���q��76�f�<��d���9�G;ŀ�+�.T���r�w�1�G�H��CȠ��tᗹNh���2�{|��r�.��1�V~gS�������v�I�H2��e�Q�tp�ꠁ{�{�b��"�����tI�!'JK�`�	�K�Q\���;��2����Bl�nZ8o�̒m���0MX�����9G��&C��֖��|�8V e��3�Ymtm�Z��{ӣ��t�V�M� ��?c㐑{�����P�!?ϡVm�����(���Q8�T�3k�K ��T������|Z��i�Ǳ2���:0�͑�����L������G	�DO�36'?�� e�u/u
��兦Sc�+�͟
�1��Շ%GE�*��+05.��� ���Eh�Jyb�{���uAd<y�_�z!:N"6����g��Ǖn�U��9�T"O1Ee����q'��g�68��>�x�6�_����h4��<s��=���7��kݳ�G�G�uG�	��;<%cmo�g�<��O"ֶ��������/�m�5= �P�P>�K[��,����X�G�y�5:�`���r=�97�Cm6��S��T��}Y����g��k)(+Fo��R)8l�%�%����3bRD��%�%u˔vyz���+�F��r> "2"�"�Td�:�Z12���7���nT����r�V��ԏ,��l),�I���tq �T'��v�'��\�����1W:R<}�<�A�CL{1E-ʤ�X�w��lᝑ6;"H9�x�b�Ա�w�7QU�	3�� �Y��NĿNib�jԫ��nU�#$�%D�i �M�����݌�;��"�T���-�EW?�Ўkb?�y%�?��ÀK��b���o1	<�5)C�H��o�8���?Iϕ�7��
R~
��z9��I\�;`�#a�"�`�_n$�S���:6u���,� ��]M+���A8��/��:dp�����-��ħ�S�5����p��3��Z[�as���_�jg�|5�#�K�Qp��;)�Z;�V�Tc1FREYA���MbP8`b��w��nE#�\_C��v�]�\ە����>��PG�	�1~B?#�K�9�Y����~~�L
bc�X�e\qi9B�uʍ���}�8Q���dl��B �j��f(�ҍ"#
��ճ!ω՜p��w�.��~�a	}$͞Җ�#|�0aV����Gg���\�7b�T�0���4�?C<���+�E�ҋ�i�VٽYZ �ur&xf����|�l9d,5�F"E�CZ��\��C����f?:5�m��mP��=����b��Iq^]��T�kFғ�JU��n�(:��mE�x"n�\����h%��X���+��v�.?��>)�VH���o4��o�L�Z&D����|u����J?Vk���d]p�'�rn�T����U!��Ke�M�Ǫ���SU�v+��%�np�{ȫU$H\|0FA9� 2��q�3��B�
}�O���Kf���h�00�ٷ�����\�0��?�V��{��>����\ҙ�hʮ�06y�$`y<�d�3���}��;��3������@�<4�`�$��xG���t ��:[�_?A�)*a��bǊ��E�fI���HxӒ�ĝjJ��L�]i���I��pfo���>��.��$bӡ�rG��/}ml(��*���@ne��1�M��7���\w�T�E�=܉ !�����K� ��-��d��8t/5 Pt�+�c��)@���u���.�%W�]
���x��W��$�2 �]8mb*��-|i�c��`K(��'A����j|�P���S���g����+tj��O �&Ig�c�(Ň��7�r�fd���Ľ0�y
��{�$#�����Ⱔ�X�ZψS{o�����������ث=*駐��$���V�/U�� V��^k����QA�r�T����W�h(H���_F���w����H$9�䏯t�R3�~������O^5����������Q��7�����p�b	v����� �%��~8+�w�>4��|�� H���m�u�� ��6x,�ܳ����_��|�@%�e^�#���^N���8�DJ��˲�U��E�r�� �o=��D)�"Bw]e�N���:np.DRH�3b2�EɚZ:�c�?�~��`�J̸�5�E��&X4�83;���l�M�2�~��Q4͖ؔ���/�^���D�L���ϻ��㸷�9G�-2<���B��Bb�_�>�s�Ң�w�E��	�u���>�&<��4�'Q�˴Z�����'��	�Fb��Si6��t�6I��^K�" �3)#�e��I��i��JV�Q�����,������.!��a[�����#=�����x{rhP�_�Cyf�>�XۆniOrC�ȱ�v�Q_
�~ �_������:�-	2� ��I1���	�>l�P=���Y�v��n�t��"�a�ܾ%��υ��̂��ց����4�ЙvJ���Jhͱ�0j֐���=����u��ݴn�c)��[�Eu����X}�z.���ط:0��c�C�/O�*K�����VX�'�=J!�0W
P8�jV)n��6���q�vj���K�>ˏo���73V����GSV�Du/.v��TY�����o��i$lX�K���uJ[a37(CԺ�m��~�[e�!0���c܅Z=�|�Ǯ��:�`�Cj_��� 	[֮	X�q*s����C�r�Bm�O�m	D����tnas��KUG��@�WGƐ��"��#C$r `vJ��sG|��%	���>����6b�<�o ��mpD2I����X}"�8��G�gFk�Y���=���1�?�fz���0��=��p�0'R�N��� M�`:��=_�c��MZ����I*��-)��@�Qwo�s���;����{�5�>�Hm��4�;:���ƒ<s�@L#��M�h�#���5V5����/%Ĵ�/٫oZ��l[��H�4f���/�W)����/�.�����(�r�:����iA�^�t�v������Mk�^���ǃ$�k�$�CI�7*ui�v#��qOQ�4#ӝ��!չē3"<��8KN���  z�>��k=��'V��I>_�Z���bʜi=M�I➫�[�"v��y����2���	�F)U]��@=������to��!��%�dSxk��r��Uq���Hfzi�\vC�O �[MY�k�f5��K:�p�l���#��J��������r�Ȓif��i�gb�p��CT��+N��S��p/!���]|\R��K�����[�|��ҝ6��)������wc��Fk�3��Of����U�^��I�2Tf�W�^,rX�no ��\0�#I�;��E[�p�󖫩u��{�����r�qH��:��(�3���6�t��t��i�/Ru� h~򳁕�Ĵu������m�4;�iG.
��"�'���k��E��®%Z
��=���T����u;ZwO�H>c�HRw��kV���)��d��38ͷ�zs����<�JP)D9�=��!;��n����<#]��e�|t����@r$��x:�7G-��d�,�!��۶:�ݭ���5�V+	���n?�#��<�(�L�d�X�{u��.?>�;;�>)#�)�X�QW���>8F���K>:qg�����?�a�羫v���ka_�m�s���CQ�����c��ٌx �R�,�x�v�k*�>�z�K<�%�������D5�� ���~_d�� _��M����bZ�3��1}S���e�ǿ9����:��Tq<�aP������>�!�$�ͥ��z���T��%��D���E�X�&BRآA I����b3�7�U�����D�� ��?��)ވgޚ�%�΅v����p���|�MA�t:��׊���͆�N�M���"Nk��b3/�㟋�����ƍ����4�\��r5Щ���\����fgS����%d7V�V/XW]w8��7�tu��r18�n�my�N�qU�#��S{#�Rm V�KiB�²�rR��~]��&;��@��uX��r"J�J�5]�D	�'���a�s&,r���=B��*�;k�������-n�z.�鬋�2W$�W���rr�f$h�p�����'R=[&)Rʓ�ǇY��I�?�*hl:Y�T{�ѻԮ3#��Cgt�̶ԼQ^,�i��ٓa��7r���<�J���!Sx7��I�o(�N8F��Y�>�5��~�XEh����_��a#	l����lu3� ���6���h���z(�XB}�է^
j7���<w�͏����&��@z�����y�,4zn�s�4]�_�.LJ���.y~*pjc;4N����j�����f���%�,�(B�.��|7�\�Q���2Gfq��deo�r02��������6<��n�E}��`[?��0c�8Ϳ��QeFJr�)�r{�iyP���M�����ak8�����]���Ku�F�񖞂�~�]���nsF~����FҼ;�+6��OP�tc8�̘jcg;�VS���*V����d�0�Ob`J�Ŷ�v%�.]���S�K�"�qAsȤ��i+_��/��;��H�?Fw]��1"爹�D�f��������iqt��"��«#�!\����<�%��`TOC�ѿoY�O%`��^B ʑs�1Q�r��l���㎮� ���8���~���A��[�), >�3�V	�,D	m%=�o���}��N��\�J`�w��s�a��uIɘB�l>��IV_�3/q��K����+�Xn������#)�J�9��M�5����= �m��n�S�={Qێ_C��X�������Bhs�}�m���Tq�x�iryTv;2f�w?#CBos��""DP~e\]I/�o8-ߘ~q��my��92E��E�񵦍'����>8"xK��:N��-���&ֻr���}������U� &D����!�R���!рpdD�I��E ݢ�yؔ��岡��Jb��sO�1�<���~T�E��7ˡ��`a-\;��x��e^����N�y��zd�$�4E�2��ޗo�CM�o[�^4�tf�g�gѬIo�p��y/�S�����Q{J�R�Qǝ�Ǩ�d_����6�����XF��ъ粕�_ruv�
D�n���cj ��g='��G�x~p���A��w^�T�U��(vg�l��8̡�cf1�>|h����D�h D'���s���"O��~��/N�m:9� Aw>�(�q �	 ����6I������Cǒ��w+���Ѱ����6YHZ���1����K!���׿ˠ��Tr�����P�IEH�q�q<�ڠ�Ы��kM�W�o��kh�o-�A¶9_|t_��Z	��2{;W�Ap�:����[�_�4W�������^�q�+U��{{����q?&�۶Z5��3�Lk��[�c�+s5��$�2)q�{��6��;���˄%��a[�� T���$���>��0?�5���O4�j|*|�}f�D,w�� ��ִp	����
'@G�C����:�h71I�� 6ع�L<?nS���LM�OM�K\��6���^�]h�,8�%.[��Y?����R��	y�����W ��;�r�	��x\�rÌO!���G���{ �/��V�cRF+�&�T�&����}_I,i���������b��Ίz׵%�>C����t�4;�N�ht��jw��ʾZ��ͻ���������?���S@t�s�\�}Tw��:]8�{ S���/��8��H���zy'���|���u%������ZQ/�#�X������g�ctӄ�&0�����ʉA���ZZ��4����n��d�5����kQ޵G�]�]�z�RQї�B���(f�G�}����Iр���T��n���Kcw7m?��f+l�	$nf|��u��1�ea�y�A��� _$J��!g����=���,;gq1_K�w6�{��y��ִ3ֹ�c��+�QtA���N;K���}�����{��yߏ,q�b	��d�^6A]��K�8|�f	X��,�̝�S���YDK�|�h�,�w�)���	5L��3#���gQL�|x���	ؗM�d�d �
/�}i�v�{��x����}�w\F-<��3 �x഑&�h�	À�a0��p��w�BS��l��{���������>��;Ã���Uo���Z�_��?��pW�A���p��,^y+L�9��i�r��IU�ސf�%|.:,@��X�`��[�MRnC9�����£��-7�\��B�/ޯۘʛ�$�%>�����+�-?����_l��Uz;�R�ٽ ��^��yH����7�B?�4(F۶���^fE�{Ky���~����-7�B]N/�v}W����&E����*��ŧ�Sz����iW>���`�Km��V��I���o�A1��4�[昻���Z�!i8M^� <����E^!}���%���6��W��|&�M��S����?f~�Y~���#V��	�Mw	���R��c�w�s~_a�����r���Ql�.C���eK�w�h���]`�*�� �/�����h�ݶ���E�rQ�w�""��x��g�M5W �*٦UZy���~�Ϳ740i՜���t^}�bu�µ_L*u���>����sU�����)�Pc\�d�N%یK�/�k����5���>x*\�1
�!�� B�{ta)��}v,ty9l�R~G&'�0fw@��0{i��C���,���n0�T���_o?q��x��ڵ$���)$�O+�^*<P'C��D2���w6�"�͡p��۫�R��ؑ7���!����O��!*�>5��q�Х�|�¸6Y!"�d�g6�<�p�����Q^K�L-�Q�ҹk�x39��c�Z�e{�.�/�%V�׃2ҝܣ�P�ݚk�
�IV^��m+(x��Pf�=�X����a7��͵�Â����ݷ��a�F�������Z�A��H����m�����Uy����2�2�6j����!����9R�'Bz��#���أ/18`}�����2��31��9���8�?��w*���}���9	8�}�=Q�Q��ע���c��j[�k���(��G���
[�Y)r̴�0>K������26S�E��bX�
m]Xz��՞�(Fo�6'��,�AQ��z���$����f��dk�R�>����<��������G�j:8)n4��������f��=h$��DT [�S�g��"<g~Jg}��7��1Cب�����l\��}�R�غ
*e��.�/"��1W|��x��0�l:{�Zo�?v�\P��${�m�LMQ�W��z�|�3@��bs��I������AX�[���V��ȻЄ����/��wQ���i	°H���/3�x/ŗ�WK�϶�M^yK���b�cS�w�B���}xv�y�5v�/��`��s�����X���d���/�^�X�W�d��\��87���7�s�d�J�|M�	�h��>�Y�o ��S�V��`����;����H��H������ˣqgG�pF�����������M%ݥ� X��Z︩���V7��E�_����E��$��K�k��7�"[��T=�|��&&;���1N]� �(��6:��D���{@q�	K_qmSڇb����(rĩ=�h<�qr,n�+>8���^�/L�n��R��r��7��+��*�E��b'��̽=L�=��l��i$ԱLp�,DA��W���'��ɴ��z���3_5ʝ�}k���@�TT�_�� ���� )��;�}W��� �0}�{^�΁�&70���-;]�b��T���~S8ފ)0c��+-Ŋ�g
�?�N�Ά��*Yabң��S�Zƥ{����U�*|c���d_|.����8Jy��D<�@�I�U�[D����ZOq'��m�����,nz���2��|�Ǔi����6񾭏o:�����d�G�턦h9L��0���0B	���Zp��塠�?�%�x����.�T��� ���i�2M%��z�j7�?~�0h��2��w��<eQP`��aͿѳ��:_/�ҝԂ�~E���k��1�@�� �f��m��1?���O�}G�}���dQ�4i�����Mz�3�B����"�?��%�"���9�d�۩��<���@A+.򌳭�����p#�¹���\Y��+G듷�1����l�c�����Yu|6�͏/Չ�( �D~j�Z~�wQ�6x�?K��~t�rS����,�-y���͂A�RNq"�N���t[F�>��GO -�$�m�yY�&�b�/����qӎ�u��\؛��[8���7��#芶QSF"߆�>��j�9���UQ�3�۱B0�u��oǷ�t�"
y�%�[��#�o��k�>�O��`�sW��|�h���;�e�~ ����ˡuPF��3���ܧ�@�n{��v5��N��`�$@Ő�[j-�a�ֳ��o������U!	�g��ꆍl�U���s�p��;'W��d�ڝ>�{^����
�9SKԿ(!8,�����O �L��PT��߹e�P���q?�Uü�r_B�63����s%�Ν�rs�|~l�X��"�ڼ�qM!֩R!.�씶�s�"5�! �V�a�����.��j�M\����Ƒ`:d��:�i�w3XRd��BCf��O�[꘭/�żMe���r�q-?�(H�����h��8N##����(@�&��xYyK�pr7J�{�Q��1��.�Y�1�A�p��ae��z/�9ɳ�w��w�ś�U:M���>�,�|����H�.��5��|v��enX������h����U磪�K�GR@g���"p�g�6��]i9eO���_��+�W.
�w��=2��1[*�}a�VIf\�U`}h�#z,a[�J	����`x�ɑ�C�"+�Ů%Eκ�s��ڍ�~
�'MY�ID�+!wKVC"�$^�����hv6�F�Ð3o�rWr]7�tH4�Q�Y2� cg�[j���~�Wlc�݇��x)���,Ba�Ѫ\��J�^b��6���F����ң��`U�S��/3���|tt�f@�W������V�,"?�TFe�vQ��t�a�����[*x��k6����9�so�#�:v����c۱;�}��e	���%��B�hp�����RP�:;��פI"Sb��~x�H+�9��ߖ�J��t_\n�� Ǆ�0�$�5�,�Ap<Ք%֜��;u�<�p�F�ߜ�n�=�L����\K��M��2��̹l1@�iͥ	�^#Mǔ��a�h�u�����j�M���#e�k�i =>]��r�B���L�T�N�cR����%/�������u��4��W��b�,���_{2,��������{ (#�\�MGS�����%�Lw#�c�ܹm�TI���Tw�m̵��og��1�QAK=G�+�uT����HH)���bv#pA��'їC#�ܓ�8R�w�\Fy�00�w>,*��)�0�jaJT�E��oB�o��Bl��r�LV$�H/X���/�R��I�}�����5bI>Y!�>��;��6Ρ�u�j�s��ܔ�.)�jo.ο?�Ѭ/��['��H���(&��)A� $���e�Ȯ�%q�C����;���ت����j�T(�ڔ����λ�����g��w�bn�g�F�BÖ_�����q_����e�Q�7�������%�l�o/���F������U[�23$X��{����$1s�x��h����}7�gٺN���8B$^+����!]��E����?1u�4����m�.@W�,X	_�V���r�V���e��Z.Lۇ
|�����e'<��]�j+^(Yt��O-C(���j%�ލA��-���'��#��͒P���_2�C}��:|�~�j����ϵaLvQ*��l� �?�����H�&������݇�plu��E�QU�����	e���`fBt1g/�VEa9�AL��L��BF�/Ԏ������]��:�����{���+&�+<���on���/i��E�V������ٿ�*) ��R��/g����$��ߪv������!�Q��
�jz8���0"+c�v����ώ(G��5i���0��C�F�*@��7+a[�7u~n��|���}xyJ��
��࿬�}"�e�ɽ�U����!�(y��gK��ӎ�\h��K�S�G�{Eʝ�B
��k5k�2׿���+�S��P�1��@����v�J�MzE��<9�%�\�������.�n·j�?�J���U\�+�*�J�j�g8`�|�����2ں��ET��h�w�)}��H���U-�����Gw��c�L��mF�Ѩ(s�G�<���Gh�������/���E���ߨ%��2],?��o�vy�����|sQ��&k��Y`�D�4E�̐������n�����ɷo\����/�&Ͽ}��51ii�'�ә���I�8) {�=���|��ʇ�[CC�&nn�A1o9���-��H=��XM�FS^�F�2��b��F���CB��ĠU��Ҙ�$�Ɉо@��	�#���v�z���z����O�aQ���4f��K��Qi��y���'<!��l�[�r��8ha�>�t����8��������땗��E�� e~j+�{]��v���q�,�#fE��͔���$�~%>[*���T	�[�&���}T`���ׄ����w��돾����6������5.^����h�~�o�w�R	��.����n�G #&�(wE��j��h �ὣ�\��˺lYr�uxK(����oW_��۞��؅'꟨��ϼ�S>ͮP�C"���[��b4[͙�z$\���������HK<>��0,���ݩ���y�/��ۚiEC.e�����Z�v���@-}y�w˗"�AW ▆ I�E0����vd��X���cBxq?5���u>3�r=,�wu�HE$ul��hH`4��S�է7��W�_��f�mZ8XU�n���a��j�7A���șrX�	F�̩T��9�o�HO�G���T4���R�ˣta�b�ٞtq����K�)��:	@y�.�o�]�U�!l���R:���u���ŠI'm���N��?�*ޭ=�ήm���
"�*{\Y��ҧ.��{��NւQ\�[u��:S;��]���E#�Ӝ�j[`�6n�K>Ǣt����H�i ����cX�I�tY'c�����]$���`�	�큲�U�F�p��L���Sb���Cf��D�:�Ѝ��[�U44Ş���ty9'�	���ph��@8����}�'�Uy5?���t�<�
�5�����K���,�!�'z�6n��C9�fx��Z<�j��5`�1�Z5��~�V�e<�D����y��"�oYq�"��G����SUj�M�[��ށ�M��v}�����@�cM-:����
q�d[��>Xr��&�����g������n쵞��i�m�a��t��8���D�k���H�I[F�!se��<���S>r��(�@;�_�>*��W"�����uMDQ3��?}�p$���D�S�j�6f�t���E}W�U
��NK��Cx�b��*]�5E��d�Z;W1�w#��Ou=�:_���v�E�������ŧ_>�j �AQ���>&k�%��w�UZ����<?��&.�-�8ڰо����������p9D_�CX!F���E�W���'v�٘��92@(���x���%ݔ�s��ifj�!�^�9϶�ʼ�EL��ĥX�	��'�̉���*�#�6�,�k�l��Uΐ��e0��SD'�%��b��z�^��R5�e��m႐9�ϳ�*��p����:ǀ�ޝ�|;;���{�o8fۭ�;�+����bI'm�l�����TG���:ۖ���'�`3�/Jm�#Z�����g*�(/�\@Ѽ�A��qw-Ax����NQ;���{�	˕���X��#�/_���� E��-�z\��W�Ur��ڦ�v�U��O���� ў�9_Ts�q/=77����\;��Aʯ~�RP%Z�k(V_�I� -�i�����$o�o=k��J���6}�d��)v���.���h/�A�5\Q�w�I�L���?�gtx+�ʵ���?|D=��1�k^FU�8�0�ev���1r�4�{�`OF7�K�V� ��.&螸�C':G��O��>���e�^u�k}p*c���@Z�\�؛f���|�@��uJ "��<0�(΢xO�2�!(���^j��ݨ���=YB����{~S�z�
�x�	EI�Ĕ-����yؿ~w�5̌"���0@
G�F�q}-1b�X8*ۦܧ��l��¥"��r�p3�x-m����-xa���]1��Q��5�9+�m޳�՚�����_��l�j3�Ͽ��t��`���7@����κzq���S=l�q݅Y?�M�.�:~���b��tB�8�N����ʏfO3�sH�}��8����f}*�q�ѕ&�a�wmWv�gK%e��zq��\����cv�t�n������"ϨaT	4���hSŻ0��gŷ�[�����h�&�	A��UAс8��M�E�I#F�l���B��\����q�>���E���@�r�[����L@19pȦr�R�H~��G�ݻ�~��#ތo�u��-���Aҝ��g��Ļ�i���n����ڴl?�����_.�ƶEO`945٫�q=��F`���'��t�ǌU?��=zߖ�^kߣ[�GG܈�^~y>`h��#qw3È���#C�,���^�P''[ȸ>vef��mtH��`��|����J�/Nd����M9Gq��'m����d����h��8~��([��F�6 P���� y�Ej���Q�.{�����j�.}��&7$;(���4��']����X�n1�|��f��~x <Ʀ��OC b�/�Y��v���9��vA2;�k���%��*,������C`��A��_N�'�!e�H�����Ǹ���	)}�6:Ջ�m�Y���)ؒM��aDc��D�''��pGf�O�ަ�t�W�G�[ ���$L�#s�Q�e���q�����/dB�&�G/�JZ�j��CI�8�Rc�Oq u�V�|�q���tJMSH5�[X������-VE���Ry@����[�s2���v���Z(�$��{�:�ߣ9�\�*κJN=7 "�y���E�vL��ʫ,��Do��X9ìk15C��7��t~����HS��W	��h�6M:�� Ξ�WMw�����s)~g�fɥ��c��O�x1�Q�,��X5al��Q�\��n��� T&��6�N
5�����2^�ۚ�zؒ�Zuޏ��j�0�~Zۗ͐!��AN�H� Ev����%ɞU�l֦�g��������0�Ev#��>�>G𭀈���ibbb�MMq�̃&�gD���Qƈt�KV	���@�'U�}�s�V��Ѕ��m[�s��(��4ޣڀv׼%���'�SJ�%~8�z�۹T+S�������6��!#����ml�tҎ��ᑡ�,K���~��:��!�E'@���d������`�0kgא���
eN�o�;-����ב��*��Q}�w��y��9&��g�򟾅�ɠ�!�m���r�Fݣ1�ge&�S�ߊ��4����J.%s�ձ�c���[���[?�c�m5mt�o�*��_[��*���0����=����V致�e�+x�|���w�9_L�??�btpEIl�J i9��!K��2x ����/_#�&.$�	��f#��q#�fJ�<�m2q4*�E����Fޝv�!G2��ځ$�]��KݎbŞ�W��G�Tyc�H<,���Z$�wI���H럿������1P+/@NOh��cL�b��)�O��A�^�}�~�3�Q,\�[�����9��"� S��P�nry�!-�u�N��XF>ڱ��7(Ť�%J���{˰(��m�AJ�A@��;���%FI�	�D�S:$�FZ��������~|�����^ǅÌ�ε�u�}�V�y�+��v�e�*Ơ�E�}���Ch�
��#��v×/=�PK�f��5��C�����[������_�������y��r��rrY��v�Jgh���)��(��ܛ��N����Y���x�|��s��/zeA���VL��6`�ڋ�^���S�t.����r��>v���]��K�'����d;LWTWe�A�#�u��ϙ�M��2��F�¾��z��7>����+�)ǒ����{��['�N0 �t,��� u'�A�)%�a�\��(7n�7�aƃ��¢ ~��ڦ�p���`!����|��  I�;.��"�|.5 �����'�����ɸ#YF�����]vE�	{�x�����]���R����{� շF1�k���YB\"�)�7hY�������1+g�iCF�ki��j��
{v|������"HxP�X9E���I֕��~x���P�{�(yP�����AF�~��4!���9at��)�ӯg"jf8IDܤՏ�s�\^]� VO���=��~a%��z��ݪ}G�&��,�	������
9�Ν��+-�r��t����{�8��d���屼��8��3�4"�G��j�K5���5��FHD}� �o}�+�$��9��8;��73;�k߀���a�)�#5�鉿���8"BII	3���5���T��O�źY>+�䮔">�C���A@�_Ι�|�A���K2��!��O.��P��+Z�O�4��D���8�ԣ$5������N��|9;7~��"���I�]���y�����Qizݖ����~6���*�yo^^l3�4�f�ٖ��4kV��ܜ�9@C/�_:�����s��lc��9�{���%�R��432�f�;v@v�+� �s�+���b$1�Hr�q��ڀ���v�O~J� ��c.�4�G#��u/����R'	��Z��Ԡ���S�6u��h���g��eВ�<��/h�R�_��������9ڻ����9��謄�y�a-��ௗ���o�+��
�hEت���-x tA<I%��`�������
�� %��}���N���yuN�Z[^�e�.c�G?���J%)m�R� ǿ,n�`l��X4ӟD�b�f\Q��G@;�F�W�4�S͓����](��dOJ��1��*a�%�"��V;��pgi����I����?bL��N`Y���fd�XA�D�Z��}�(w졜�#�	,;��dr^��F]�,�7 0rvG&	��p/���F��V\�YNsk2�� ��s�9"K��L�4Do��Wc��������r��p5��,�:~@s�㲑f9C��c���Q�j$�w��4��%bJ�О����W��>'?�1���p�N�q>ܕ��x��{Yn%�-#�}����Q�rni���j|Vdu=�XU�-�#�b�+`@�T 7��z�u�% ��~$}�܌��"�����&�C����*E�x~�uo�{�ξީ���6]e�W���Y���]A�8}Ӊq��6Ru�mp��[d���8� �pM!w���ru��"v��7��k��Vn"�}���]h�x��t�������^��B��p�{�c�
%�9���i�����qiI׏0!����Z�g��q��~Qm�a�6� �h�aq��0��%a�kv��4���4*��:/�[ovS\	̾�)߮a��0�Э�H:G��d0W�[��T��m���[G�kNNs�((`<���l�3b,�E^��3�*Q� JW�=�����U4c��.�!����CmI�r���{���d�P��O]V�[껾�3 kuM���ՕZ�`�=��'��'h�v����A~�@z�k@=�`������j�� ��<|����8����B�������b�`r�:9��,g���	#�z�J�ܥ�M�_U��+���&��8�U.-"	�E'&���L���� K.�?,?s5����^H�V@Q]�M0Q��#S�sR�Q�����plЉ����s�b-E�X~įn�НJ#������<]?��4�"�/���Ze��H��!4m���������L��0]����B]�ziw�gJ9����ej�S�pp	~@��j�X�sm�!n,����N૾��rX�A�n��F!�I���:�R�K��'�y՟����b�4|���os�q�o-���� �z4��۲8s���ܿ�� ����q�w����� ����A6����׹Xx-;���|��[��,܋��Y���G	�o��ݩ����qZϰO��{�Ø����|�ކ�J���ͫ��1 ػ�Y�w�j`$��1��[X��0&FXc���^�q�\?q�X
�����wB_TS���(��Dt|�V�'�|~�!�V� ʵIe�w��X��)�L=�͖W�����@̥�h���eN4<'� E� ���#�#Y�y��Qz>
sI�Al�����<�����y��+-�Vʯ�3(_��+~g.������.:�t��;��0�p��k���ay�"�,����
��|�G��.���˔ʖ�l���T���Rm����o(4g�jT譮��?����MzYUd0��>�|ou��vDY��D�2�*��TF-%9�)ӳ����O/�=?ߨ�	�ݛI��)�{�TE��"�wJh�+��@S_���e�;ӥă$��<�﹞U`|�J���k�P�QGo~�����U�S��&F�o;�aK�gFqZ�v�# O�	���O��8��RT�y��:PC<q�(�C��9Q��ݶ��`����?��9���f4"�/;�6J��|�.���i�e(�vG�.+���f��#��D�=H�?���������3AX	2�Kן?�G��bG%Hާ� UɁ�^�nr��H��r|7����N�<���i�6�ܒ���f ���t�Rz=�Ȟ��v5���.E����f<<�P[���2,��swH��*)iQ��{B?
��)���![�Y� SeT�Oݙ�l���r��+���Q������$J�q�ڣ<\:`��ls��"�,UXf�fURb��V����e1��P�,gP��L-��v�,2�G>Z�~T?���W� 
��s�>V���P�Z��c��lS?�4 &�\���n+���|O���d�����aY�� �Mq)��^/~�,	�h�v_��J�3�uA������7w"�:�J����@F�l�fh�xz_���P执�A�ֱ`Z��A�ꢠ�;|g�ǋ��t"3��ߛNh���L���cs����݀E�媶��� ��a���7/��=8��#J�o�������F�^�� � �۶e����� YYZ4ܼh���a�p��nv���a҃�p���Vq�P��%μ�	�/M,B/�-"�pJ�r�&1[���r-,�,�v�b�d]1�݊�b��Qj��T��B��q~	k��������C�۵�W�E�]c�]��<�]�Tr��Ę6�D�M�$*�J�ޜ�?��"I���}�u��@�y����O�
|��y�v����a)֥ff�S:�����i����:�u��:�-ZFQy�2(��ج�*a�`2�s\�8�-��-߬L����ba�����9I����P%i�:b�#��"��IL(�#�&]�{!㯶>��dt�\�㙵��
Sf��X��\]= �YB�k��U5���R��/r��[Xt��vy~	>!j���bG�K]��e�C5xy�n[�4�����w%/�v.pkZ���Z�g��Z@����Y����0��#�/�m�5�{�c���U����� �ہ���q�bŴ!�Cip�ZA����6+�6�.�1�n�=����o2����5�&$X��O)�r��[�Rx�2��|=��#�V�䘃�~Mn�?��f��F$ �B�c�
+*�Sd�U�1/�F^��A��U�Y��sob�k^%to����\�]O���6��^j���r�ݖ
�}-���O�Q:�u	�r?�
��M��iC9/�+�^��L�<Ġ��Q�(9���jO~�B%�k�4�5���SpFkT���[���bPp�ĈZK�����l�,ș!�+�B�� ��*;e&�S8����p��rY��;�	���P��hLtt�����Yה������b��Ww�9I�5A�>!�Js���)'/&zZ�%���kg �sz�]�fjZV�\�'������އzl%ᢙ&.��[\t�o9���e�t�a$���P�(:��WQ�\s)0��άc��0N���1��ೞ�S���;B�շ�9d6}���U��������x��<�X��r����c�s�iGۉ�'�����л�YM��1����Y�D&��B'�C �o�5`ɻ6!���ǁD&��{2���
�\��e.Ҥ�D�^h�����v�f�T��w9QN��1i�}����;ӏ����&�"֙�+OU�x����&7 �����.��X�ו��:���N�������&:�m�=6�������b�"Ù�>1(UCG���n�q��f��mg���z��`��!��&���^^_�$7'<WLv]�n����� ��6@�Rk����-��3�/_��"q+ -N��!S:@˿���	��=VVI�p\
;4�|���y����6�ѿa�� ����R��^�HG���X��C����x�%)/L�"w�OiH��<Y���Ԯ�	Nk>��xx�p�~і����^.k>�O�um��w�ڜQL�yRt��2��}G����.Q�Ϯ�~���g�umN���+�r���8b�+3��w��(�Z�����eb멅��85yd���]p@��M�dtf�c��.�p���/�m܄,�<��>H �W�RD�,��]��6��d!���Ò���ΙJ�S�O���_�o�!6�y�[�5��/i��e�m}t�YH��#F�8��Qa��Z��SN<�0u�r�r�Q�AF�K��i3�3�N:s�.-�b`��-��Wl�bw�헞�Vί��b�X(A����ǳ�n��N�.� �@,�vG}N ����=w��t(�r�� ��n0S��T)���J���d>I��1<A�X���8F�Q�����D�\{,0���L>�c��^Y���3���yUĴرb��Y׈��	��X�U1��[�8�ق(��
������1/�ۉ�%!֥k!3��Dn�+�����D΀m#H ������*&Q�RŐs�F�껓Ʋ����F����Kˮ�I�����uͤ�_> =5Ӯq�|2P���@���ak9��כ��]�;X֗�1��
m�����	�TP��)"h5�?���EJo*Hb���n�|�*[$仨;��
��?���Qad(��(A��0��0���e��]��)믗Iӎ�t�����Ut�����z$4��)�ʛX�:qp����ӌ�s��Gl��ʰ���#�85��h�e'B������*50�4k���o#�+��H�
��Q#!�����_(C�a��L )�M�����!~%N�XꌿO�*Ղ��ܗr<�����{����I���?��[�qr
��4T���G'�q"�:I�x�!ͪMI'�:�#��2B]���4��g�V��U�*����P�(p5�I�Of�Z\���r��`���a�]Q�y�w�1��Jd��wx����{~�1@���TY�Z^I�#G'J�~Jb���������m�1�I��$hjH''��S��N��Sɸ����R9_�7���c��=Њ�Q�<��.���Ć���D��NX���������q�bx���n�Sz�;�ZfջS�D��}��BP�2�ķ�%�&�t(\/�괮[�t��P3djeC���ҩ�y��gg!x[�y9���9WRf_��4t�^c"u?2:���#{�׾�q�q�4������ɺ��s��o�A���1�j1f�e����d	g1��9�z��!edyJ�X.t��4w;�)�p>jX���Q�������إ���w��s(73*�bU~�CϤ]D����#)uI9G��#�(�Սb&�C��C�߸�ê�؀�v�sI��MD�\9� ɬ�"��?���}��qص����eOE�&X�#�?���˞}��ZU��As~!Γ��;]���Խfk��)�=$_���I~F��C%��~(�/>���17��YV�Z��id��$�q�^�Z���}�#R��z�g!�QͰ�<��iC��[(x�s��㘭�B��;�<�z���2B���L�$m)���j)�Jf�Վ��ǀh�p��[a410:;~��#0��'(c���RJ��������w��<�U(+�˧s����!��HnZ�VD���Ed~q.W;K�M�T}Q,���������v��;����bU�X��l�b�	��Cο�X_��%�L��;>r�Y^\<�$��op���?��eR�H��v�X�?�`Pph%@7��s��E}3a�iH ��|��(�1}nҍiv�!���d����;�\�~Oi�J�na��I�h��7��i �!vy���^���ލ�r5�T����\q@0��] @�^M�W�J�U^�H��쥺Eb��:��Ȅ�~��O�ƃ���^��5��L��S$I��у�>�*��kT-�~��-"\\���D����ːbGs}���ǉ'ňyD���	 ��b���X�2Cb��9�"��_K%�{�<���C_ �T��!U��I���ǆ#��?�2J�)����k�J���	����"��)V=���mj�~(6�Eu���� DH�L�x �����w3��o�p�<*/i����T��\%�Fڅ��5��U\*eٯIX�~�yIݏ���s������������{5`�l*9��
�,o ��v���od�������r(�����?�A1zk�7>gDHOh�wQ����p{� �r�SfgGeDx��*P��Up;�^��^�V�]3�و�rv�?�f�L��9nK96t�Z�,0��oMr��Ƿ��Qd	���H'��%43V�DE���ys��0����$&��E���E����~�q�1�W���L�|���E%!�%��J��ְ�S���5�C�=��aM�4(~#��-��'��[���+�[�����6m� �����D,���ﱸG�0.�+�-q7��q�olb��rtݡ\+y���7��y�#�����q��'�����Ȁc܏�B}7~u�8n�\4qbA����-+�x���N��i�Mv!���La����ªS4�iYq=���J�4���I �FdKd�}!��c3����������Y�A�����Rb6�T�\i�b������ `�R�ַ��[E���)w&[;�� ���Q?�p�9�����Գ����_�=�������ZFS>F=�G0�8��\/Sӄjq;-����3�r"����gǳc���Q_)wv��Y�jm���p�����(��z
"�l9�!Q/�~n�c���.&�:�`�d��y����x��4�fWRN�}6Gַor<~��6�*��x�j0p]/?ev����C�<�'�8�V�A'�:������j�����;�!�����_������!�Xҕ�g�]t!��4Ag�mO�����Cli��8Խ¢�llV�G����$�����P���yt�d�yZ�HM���k�s�ojٞ�j7�z�8��_�uޓJ��&��[�ˬq" ��G����.�'%� B�ZQ���с-�Ah�\�$,I$j��5P�:y�8�pȥ2�,��r�^�f	 �W������4�^���o�ƒa�&����5[l�HߤV]�S2z��;�?�E��72��YP��n'NR�	�|���Y &1�g�`�����|̏��K�ș�H��| �Z�jv���b�g�q<�J�	1�����8ET̿�#)o��b,Zwu��',����d���mo&��R ����̧5L�5,�����?㞗���_V抠#i��"�ϑWbe[��$�s�?Ǯp��R�7!��LH�-K9D�Xd�m>=+���ƿ��\@�>�ڦK�'=@h�V��M6A�p �"���H��4�x�D�y�=
���D�'��u��*����(�R���p.�Q}x���>@�Д��Al�l=\�3����`)����G+~�j���ɿ�J��t�R)_v�,�4�n�Z�~ERg�to<7��a3���B+��6%�{��$�*W��K��Uz�#�^\���3���ґ]�"�E*	͘;����t�>�^��Jy�P&�]��������]�����<��9�� ��� �Z4��\�0u�|���)�P����Mѧ1��=죗���_;�݆7�^�Q�E�jP:�<��a]v:p�r_T� 5X������R�=[��uUÖ��6\r�K+�;T��
��/�ؐK�pj���q
�/�2{��D���$P�����L��LN#���b9@©gW�譹c�y��8�ɲ5�jb���<�Q�撸�%��p�� $�>3�@��]h���yi
��B
DA7,S_�,e�ȀVZ��gh���rF�̡�uщ��%����ݣ#��ZJ3"*����66V�1CdZ���Յ�U'��odte/U�E5'��S�9� �ac��gimE��f�zn���N�q�]XH�"+�*�D;�R��*Pmq���1�����+_ͭf�r����9��Y)�R�wÔ�ؖt�� ������`���j܄ޖ؈; B��`��:�i^�q�O��OT��5%���s�W��G駲� �O��v�Nai�0-U���7P`]�AS�A�S�O,Eu�e���-�	�2�iK�Z�IGiő�3<�1���v�x&`�,ќ:�3���c9�_��)�����S2��  |N	߇�� Jڨ���D���Wvn����H�$���>Ǩ��Ƭ�ٖx��論;��ܦF��g*w�z�#Y�L�5|��������e4�et�U��U�����!�'�R޻��u��.z�,%<s�]ˉ%���舁�J�<�8��,�������cAY(��,�~(�1�E�P������56�"��ϥ��������CR�]��x��-�Q�$�Pҗ�����7��S��|��\��O.?Ha�������ko���Ɍ*�ɬ�M�;�:��|��s�c����l�B`����Y�T f���{��T�����*�'3�*A�71�?ZHh�����a�3:�b��J�OU
�G��#���w#����ەS��:�_�#��/f0B���=�B�A�����h ��D;ƌ�NN,2�]�y�������N��$�z�2����U�!��F����b�dL��K��Jф�MϮ,z9�s?���
���dY:&à��P!������ڈh���)m�uh�I;80�Z��`� Al4���]�C��a$Q(H�(���g�j��3��o�2Kش����o�T1(	)�ۊ�(CY!�v4N�����s�Z�a���9�ẁ#y6��3s�.�z���*�3��20����D-XyB�����G�76�qE)@iy��8��8C�P�sE	��!��A�8XdA�Mj���:���aЖI�F,�PM�ޔ�9���ҵ�Kz�����/���d
�N�?������珗!��
���#J��_������q��o��~de
��>t5kGs$��Vjo�k ��Jd���ƣ�,뛁��~�M%(��rJ8�X1�.v��c�����c����sCr�ML�RY�N���׼��B�����Kѽ�����,}�� Z�S;����pQ�J�6F>)�p��?v@�wW'�	,����C_�zzz1�Ro������q�%�e����0Ҙl���c��X��F]ʰ���|V��xi*aC�Lq��{|����xjآ�i���(+P�{sл "A�gMFx^�xMF�x����x���Hf��$�JY�(����%v	��a'��AI*�U�<cy���VL	���gfe�51Ɂ1�muÏ�«�����`N��K�^���UF���d����k ���D��Ś��H��A���|���.Bp2AS ��Vnt��p�a���_��ŕ���*Mn�)��U�Pr�h��۷�C^�-���Na��Ӄj1kx�bkm}�ǮYD�H�z�al�&���Ԫr9�*���}^qw7V}�*�
�ʦ�J���b�&�Y��KGL�`,T7���Q��
؅X�*ϣ٧�"і�@+��ߙ�9�1 �B1+ˊ'kͫu��O^�H�ǓGn'uzg��P\���(܆U�|k�!��ɢW���}�i/���\�*�+��tD���W��k�V\\O�l��pN�6����M���3
n�#��S�O4��U�
GF2?UH�bA����_1���g[b�i�e�B���r��ȫ�{di!��k�vժ��!jp.bMD�&�z���B#niXDH_��9R�'�[3k�H�{,�y,Թ벟�	�4;�#�1E\�UNçJBwk&_^^�kⰲ��M��~��a�O��,��������7/�}o&`�.�P�P�����0��Ĝu�]?p�M�D|j{ij���0Z� p(4���̌�R��O4��C�>|ȻJ������2yb�2���ڝ7r�9<�>oks��4��̏/�46��y�A�����'}P� ��3��w�[����d����9X4�������G�p�>;"��c�t�.����'7�������'��9RP։���=?,���^�4ާԉk�2���+K��З���,�����2���g �D	S�������$�<J�XXY������_�Y� ٰMG}xpՐ�(�p���{�sz2��L�o	w�טy�B��}�ׄ���˷��k�y���zN�%<������n&ț/zps5�� z ��T�۞�����t�'\Zqx�/�da�.j�>̋���j����!~�����"!))���#Dct�������0�����''�oֽ����B��6OD\�n��r|!�!�f��<��8��'���De��+b�|w��jP�݀�[|!�����9շg��o/@�zi����"�C�֮g5�W� �������t�5$�mO%�7��ٟ�u?�T3���j���x���䓆�;��Kl]�+G^̰�(I�/k<4�$��kj��7o2�N"xFܚ�Wx�,���Y�x渷�!���k��@�,�X���w��	�]�/��xC� c�� �rs ��-��]�V$tp�2ċ���2v�3ο[��1$�hD��x,�.�����{���sj�h���~nڭ��4"�;��M�.jh3��A~�8V�:"��0��'��ڨ7,��=�e���ķ����p��t]�oN�%1I�(�?<�Wc0O�+�(~f)V]�>k�n}��mq�# ���̈��*P�h�0 n�l�	�ytU��Z�;�r����f���b����U�Y��]��̷R��e��:T��|�p0��S!�f�n�Y��1J�n��;�|24�y�6�U��c�y�5P�|+s��d.�;�auV����o�3&4���Û��+�:�	y��Ps��К��2չ�]��DYlZ��c�8��p��$���	�<�'�����m��,q��7Q	\�Y����nܥ����B�bM��[I�E0��А�5��f��T��1�ܶ'�25�7{w�!I\%+L'B�uQ!��g=15a�Z@��մ-
�@�R�,�o����ON���W#,˘��r�4Ù����jas}5��_h���Ŕث�:������o��q��WR�zn��~�jSYO~�v�$O�	0 ��?�������wB����t�͖3��@�hG߿;HU���Z"� �}����j7�gO��)m� <`.^p��
��0K2�zr����z�.O" �X�a�$t}>J<��Rg( �ц?2�8n�{����k �z	��&�Tp�-z��4�ɺ.`2ſNZ���Q���5���	�3:4�ε4e{U�Z���]��?��U{�����ƨ����r��8���F'ʦ���?&��U�%�^�)�l�(M֏�l�RzE
�Rt!��i�4��F��}�:���g�����3�[���*?8D&U��
��	���P����{^pieI�,_���bG%����������*W5򤴇��%e`�����bk�
x��]���ԕ�}Ο�,�C��g��h�Y�9<�ì��E�y�u�%���_ɹԙ�T)z��~`4l��5;��Mk�����KBL�$
�F�:�tٓ� �����Q� ��ҏ�`�=�rM��O~GvL�0�h����"�,Iv�U��Rn%H�4}X@���}_7��׶O؈��NQ3z��^re��FUד�;g���.a�dI��U�-��$3��$��#Ԕ>s1jr`�("س�f��ӭ���^��Z�ԩ�klǕ�{,�"�K-�E]%��Ts��w>c�GK�/�o�hP�X?I���$�g[Q@���n��r�X:��t�*�89�P��F
�C���ۇ#��x�hW^����Κ�u���S��Ks׹�����v�pٱH�Kӕ�F/yS�n��2�a�ۆZ�F��Em�b%����I\(���)p�}~���f�êo�ݾܦY �>�x�u��G���:ꑯ���P����sJY/~:�PUlT�e�rhL��x�[��q�|�z_g�_�.�?.����
D�6[�]�'�d"4,�Cc�+Y"e�#\?~�)����3�r������n��>�լԇz2+d_�3W͞�(��rD��c���"aw+�ی>���+�-�(ݲ���}��3ϟ'�:xۗ�"���Յd@�;v�L[f�����&�������H����i�;8 ��'4hI�p���|�#Tc�������b����Zlؒ��bU~��L���esa�-~RGO�~T��[�=�[;�4n��P�T.��-�ծ�Ӟ-e����D�,z=���HI0�a�1�u6Kp�p2�uI�3w]��[�IL�5�#��<�ҥ��+6lQ����y/x��o�<&�,:]k��qu�f1\ڥ���Q�ӯs)�����3�o"�K��F�j�U��b"�X�4��~�r��щ�iK|�z{����?��̚�Jl����}�U������@��z�rH(:�׷+�r�����X��kS��א„�T��
�j�4��W���-.��1/�>0~&�}�HE�x�,�a��Y���ON���(Fx����gse*3L�0���N��Ջ���DM�[���`����ẖ�W��\Oŋ�$��?�oy�{Di#�I�X��RBć痾[d{M��7�!��Ԥ�O��t�@���ח�����M R{��x�N?Q�M�:��Er[��0$��|�!	�X�
�,�6K11��PÂo(�)u~{3�PwO=�A$���`y)!�����E��y�)1e��ԯ!���n-��~��2�R<�$�%w�r���Z<xNr��؄�_}<�ZKM����Nyh���s�'éA�Q���$���x�%Aj�t�N�i��;���m�\J��9y�8�UX�t|�'���4��I���x��}�ç����q�'y�]Tj����j��.<�^,��	�ړm���?�l��2YCG� �3���x��7l�Mʷ�Q�&N�!�n�΁{y��+�<�X����}�x�I�ė��p�<M�?��2���H,�G�%�D��[5�96}���l�iv������M�~3�x8]4�1m�Pnf�,56B%j�R
�%�vb�e����COOK�O�'3:���2�b���?��������a>1�E�&B�^h~��EJy�d���u9j!ot<U��rJd||*�숤-ƴ�+�.�~�9����Sw�k�y��y�K����G�%��Q�� B��:&x� �b����\����W<J�cj�e$�2�DD�S�aiN.R����_%c�I�)f���36E�wV]�'D}k�M�J���6[�@�9|8W͎�J�GݟK�=fP��W̗-]�b�LG?�!���\���l�}g1k9�����x�3 �I�l�����?��y��f���$�U�o�;!���ש�����3��0�+�SY���.ޞ�hpX|F��K�l�����F�AXA=��||�cV�Z�" uM�yR�55���N�&r��CQ7���s�
0L�mI屳���$Xz����aG�F�7�[��_�qUG=�^���)z@�UzBt�i(,[Oi�M�����{EW���g-�?�~�hx���w�վ���� �mk�urL�S����~��.-n�!0͚#���:B�"��9�A���VE�g��k-O�!�2��q�ڹ�A��y��{ħ�S�h���y?��(���R�;1	�t���"s���54ZU�,ltFD�.�k�y�;�bO.�LI�@�#"*XP�L=����g�ps��F����:�:g������OjF�Fr_�ޖ�/'������C����uޢ~��XP���N��*A
���Nl��+���������?k(�����n��(�[Ԅ����j:�gN�:�M4���~޶����Kܢ�p��L�<fu��Sٰ��՘A\�֑q��H�&�ȇ[��zʍ��,�I���u�3�:�����qQ��~��+*B��υ��mЊ����Q�k1_��]��~yEZ6
Y�_��T�@U�||zE�$2U���(�۶��u�a�i}-�Yg_{�p�64v/��������y�2i�?��]���X��e<^�;��������ߨUZ��TlX�U�R!�����v7�ݥ�d��%��wv�y�f�Z����jGG���	U�߼�=�A���
�ur�$�\��_��/?�ou������d�k ��3��0��_<؍����,�z ���yЙ��i�: }��<#���RRh?�?��w/>��Z˼�CO�#(:���}pu������6�����ĜJ���Wra/.܃�7i�{�
�y�%`w�W���Ґ7�+�A��}�Ń%�#���
Pe,���z.�ܙ���f�{��	Nb��j�Z������Zd3�4��]%���:�I��G�/0f�K��D�gC#?�0;�DԷ�7�Y�n��8^7E�}Ȑ�C�7����+:�5{����������ga�C�$ ��NّJ��_�H��`�g��&�>G��@׽,��]�ԩ'��N�:콳��"�^?m�
>�o��\�GF��q�u��*�#gp���JQ�Ó툌^����T��b��ABt8�n�s�,YrFf#*��M���з>?7T���W�ު{�,�w@�n�}���oA�=K��j�� 3�����8X6��z��� �5'� �Fz�сX��,Ѳ?[;�1�����Z1�7����2��_+���v��S��F�����NJ���y�T(�V� S��.e�?doVT#N��~��%�d����_�B8�tƱ��=:����x܉��l��}۬^�����L��,��7��EiA��]��kB���@���l���t�6�o"U�'xpZ)�� �񼽀�{x}������(:1�;q^I���<-3�ۆgx_+�)#��/�� #-��ދ�_?�vn�ͷ%��N塗�;s���e��Q�&r�>k���Gޒ3%��ۦ���	Uc^����Y�xc�1ѻ�$5�)����0�#v-P�i)�E]�tWOg���JĲ�<�;���P�]��Pr۪.;���2�ik�Z����M�g)E�����r>��@#�d邡���iU�}5�{��'����ib��՜���R\"WS?��ů��@��ή�Ȼ���e#]���Ӕb��S^8��L>�G���%�}�8�4��{1	�K�i�
�Φ%w�����J�[��F���%�����_�CGAB��t�;P������t�a��V9)���K�F�/��� "�i�7+�`2� ֵ)	i��w�P��h)ds8q@�K���v�&<̆��R�r����<=O�>���t���*�����;���8�^1��888�5��Z�?�`��,���#��޳��6�鐼��g�83�Ы��:����=�Q2�J�B��c�L�T��F&���.�����d���TD��7�?���LSO�qxi��%������B6��h������hx�M��o�C�燶(���P"��}��W�T����+��C�OAAe��s��<�)$0h3x_oO�A�H��z_�Ұ���O�!>���
~"w���E��?�������~�0��O�aλb���D���[�K�,"|�~�u��K�
�� ���8z��������Ub��;��L�%G6����\�!��I5��7���;GM3���]R ��ѻS�W�}f�5q�l�T��"�V�ćVȔ%�
�߉�����JX嶹�϶�|�A񗠛�G�U�
��&���cѥW,���AP<���$>dbM�U��Koa/��}�����X�v�
�{m���W%lt���
Ɠ0���[pއ~~����g2;z��=fո��y���;L��k����M�,'!J��	�_��� ?{y��UxۜIX����w:�*��jv��9]]EfI1Tď*�?>�m�����~���|��	IO�l�&N|�'��Cm�m������,��>p���B1-GD��+LL�5l�u�����{�UU��Z9u684�'�N)��䶟�،4��vɶ����3��Tfj�8z9��gWOO�H|#��c��6�܎��Nk��#aH�J_�˝�Fm�'hal2C��&��ق�ſ46F�#0M����O�U�e�WWG�x�,��?<}e@T]�6J)R��"�H���H�4���Hא��1�HJJ����w��y��af�Y{���]���ߪl����l�;�t�Gś&������-�c�N���x]����q��Cӽx���mDBmi��wP'�3��~#���6�y��[[B�o7
j�K)l�
�p$+j9Ҵ��	l2�E�+#ӥ,�;�p�|�Y����Osk���{*�knj������uV��X%���EPF?dï���a�nڷ�4���*��lB�p�(��]Ycss�BO7�>s����AF1�Y5�������9HJ��ճj''�`S�5w�y���ŋ���T�����������i���S)�ٜ���vG����_Ϝʴ�m�,R>�~3���I��G�wW(&'e���a��4L7�"��{D�#*;�
P��=kN<���1�gM'��J��Qĵ�la�: ��!�*z��P���~A�bs��g�/>6���l��`�(��������
_MQ �#�2���?ufo/FlD��jDq̟�K�q};���gR96e	�&����c�f<>����9���j1�bdAhqtUW��xW[���y�,��P萷ȏ���Vꠘ�m&�oϐ,��:s����k�����k :����O���Ḱ�%i��Ҽ9ӥ�&��!����u�#n�Y��&W)��0�8��Al*�;9&xQ�֪B�E2X��g�Uq���9����@��� �=��B���jz���7��O��`�= ;1W��H��#_sX���"V%�aNfL�[\^�����I �2�K�����o�~AK�W���UY#�	�岥�o#� �G�kVR_����(�6�o.++��'��hOB�l k���V���E�Y/�Ë,�:&mк�|�hA[����z�^���ۘZ"N�.r���b�<�`i�3�F��\�=8�q�vbL�H���/�yMm��Cosa�֓���G�)ҽr-��BV����=�p�	�d�	�)k�����38����).���Q[�ÿp��M�1z�$��b\�<����8ۄ��BnH�n�1ϧ��0 (Z��o�x	�5�G��^ONOK0����MM�����LWQ~��WXOO���H����'��}�Կ�Y+��a+ӱ�wS��s��(�]�aN�jg�p^e̸ ��<<a�<f�:>�=���E�>h���$ri?����/H�XtΐM��]������=�M�X���+B����B�06P.Ç�*�%*����������Z���2��5{�[AC�?�!�5{�m=�*J�[*��r`-}����sBw)����1�v�����d�����闱���w~���Xt�	>F�H���C��#�������"��f�ySnz=׼D�E���Y��!�P��kb��ȝᣮ6~�'n��gR�t�B-��"��C�T�|YU0% �<�������'�����Bf��O��)#��������^�ә{;�~�|�j;��,�W�|L)��J�vA�$r��3�$d�Zu�{�w��F��_���`{{���Κ�k>� �/����C	l
��(4�X
��ۋ%m��$�o�-1	I����|I��נW�v@�@�ŗ5_y.>�9�����2@5�c���J��Q�.�*�t;0Ss�<�1۶�h9o]�R��*NA].��-���VP�K��7β*����e5�b[�(��^�S�JxK��
�?��Dz���@z�@3����]&C�mt����� �+�/���팀�X�J�1���z�y��r�P >@S�7	�}=�6P@k�R�E�����M��{��G\'� f1��ص�T�Q6�*��_	i�����,�U���}��u��|��{;+N�Emx̱`�'m|�
�� ��?�.���0&/[�D,�<6:꟞NE�%J��m\�� � ��PE;�0Sl
��+��':#�`S3d�WgFI����P�T8R7:f��������V|���]�a��l���/*�O(�#5"@܍�K�0a��F��[�*Ro����%u6�5��a3r���Sw�l_��<=�ˉ	���
J�����j���~�.B�5�p��g!>pʠ�m:\�
���X�i�*;�ؗ���Č���э@/������2l��I�d�d�W0�i��KG����c+��}d��φ���FK��,]�:��Wlgw�pP�I<�?���'n����)���6!�zG4�A�����m�cJ탄��3E|�z�����BU�c�l�Y������Px����_m���zlp�w<��S�T%f�Df�?)�Z�5�o>����vx����Lݜ�٘l~n�{P�����P*�T5Fh5���S,*�_��$P��>�k�n�!M ���o(�Q��)�$�
��ΐ\�fI���|í�jS
�b��4W�g%`Q�����fUE�Kdr�[��*ΫL�=)�?�o�����x�"
9L���PkN׾Ԩ�Xk|�ʠω��Ə?��M$���]��$5��M�6A����Z�Pq|ͣ�-{r(+C�F\�Sk`�ǲ�X&s���2G~���l�"�w�ާw~oq��8��#&��f�;��f�W�s#r̼����t�|�H�j����_�h�R�W���"��!�.�E-�e��*�B���@���ou��o��[��ei�g	�@R��F��3�($��ջ���)M}óm��w��P䞌�`�Ȟ��������Y��-�2��EO�\��`�A�����B}�II~��80B7�T��h�T��R�i�Gt$��W�"Ǵ�Ϟݴͫ�D�-I��<J�v�W�:�a�`e3�N	���Ģ~�FKc��C�za��m�,�2�tM䔄��%,c�n�s�>ȡZ	U�q�V����|��_�R�4n3����}�7${CV�s�ӈ�d�߇�*?�_e���RӶe*v>���7V�㥍��pp�Q�i�̗���if>

Z�;ܙE�7����
�[��E�.���Q 
a������Xxsc,�a��A��b�?¯��{��z�bL���~���x��8�W��޶�R��n-wV�n��^ً�W�����ѽ
�[�2��^����yI{���)M�����o��O7����WY�-���e�p\^���[���x�L�a�..�57I�p�2���l������N����m����**�;��QL�����qQ�+M��T�<�h�$��!=�vO�un��Պ�B�9zjU� ���jt�TLgX�;���6����R��3���6��)_�$�_�����ωq��A����r$�Կ��'��Na�ެ�8A�AoO�C�x�B���Z4Y�ѧ���[Շ쀃y����kU8�QiHP܎w���'��i�-7��~Z�b��,���:ڡ[h[`�ڌ�������0�4y/�V�\�Z����by��ԟ���$Ȣ�/o�DD���(QD�~-���n���6�.�
qh��P����M6���	��[�to����p�o�X�����c��.�M=��%�A"�Y��$��;OR{��#�<'C"������^���Ŵ�̆�=A�}�dx��z��Jj͟QHړ!�,W��Z8GO5, =;hw�i�l��H3 ��d�9i��'9�������䃞H��i@��ݞ��k����t6+ȝ7
U��{sa$z���^�0�Y0�K`��=EIL7/&sc� C���a&�,:r���Di˙�$�5��ɜ��A���Py��ЇuA�(�Vڈl_gF�B 8�p=^�<�����ٚj��/	A?��0Np�n��q��2&��?����ي�n�Jا�\c_Km������ov�=�gǕ�bݎ�!=�b��ʻP��������$�sv����&L��V����'�<���0�/;�bFNxb#�|ߺlGę1�>�^���
�.K/LUF��Y��ʿ@3�����5��i�Y�J�����Kޭ��0�Ef|�|5Q��[�q؞m�y������1Q��'�o�3�ߙ=���Qcr��Hq	=���q�G�ҵ�����xV%"-&��?�_*?e\L识/�{2�͏�Ȣ��>ͽp_T���ff�b+�����W7վ����@6l8n�����Kᓽ�wF�ø}��H\�l�������1'9Lԕ��Y� '�y���W?R}nG��6;y��-'�R����'�}�Z8�q�W�=���3]p�pܹފ̠2�7�V7�Oj���5��35B���w�p�0e�v�ԥ�]�v)�M���D�i�|S���Y���M���:�A�w�F�1��Ԡ��u�`k��s��c�]H�Ha]B'��n �4���m�����l�E���y�{w����r�9�氟c�4��R��3�v �G��ոt�q����+-�/��K#S�KUU��a{fO�0�$�.�]���5z�h4�{S���L��Nɐ����oٟup�`���~�+^i��V̎Bp�Y����z֭���p�<�Ld�>$�UQ4dP�ϩ�����ba>�4������H$h<�������%���8�;�� ����~�(�������J�T��alK-:�G�si��Mk�'W0�4���7�^��O��>{g("ctxnM��-����+�aSA��º�2�B�}����y_���G��f�@�]�-]�|���Jܱ�,hm�~� ��RÃ��S���c�@w?%��j��9	��U���l��:�ʙ0��^޳�=�/KG]��o�V�4�O[}&�& A�O��J�!��	��w�"п�!;&�d v�c9�{<�p��wn�级CH��Q�Z��_�9��t�?��& ?��Cb���K�Z�� ����;7�� �c-�qA_/=\>^���"q8m�l����e�Ƭ!�$��>�W7'��a��i�P���`�+(Twlq
d�+���žc�9�U�/e� �M�$�8������L�/w�LfK�z ����0�;ߛ�ԽNN�6c�i(��ڨV�[@W����v�C:��v`��o�W0%-����F��R�M�� �<��v)�e�p�1��e�8�%��bl8dJ}R*R"�젩�}=͟^�g���#k2.�����t;����*��U��lg�cl�RĂ��\I�~��1�oW��,��
�M�����D|�&�qI�����ǲ�oQn�.�T(*�A��Bx��#�M	��l���.�)7�&��1ql��pO-w"F#Z	���=?�{�v[��-��w�������o��gQ�}	���CU8��0�ԨH�i�����*؋<7��N�p�h�GW����"K�ھ�H����\��{8�~7��P1�/�|3�C�d��Vvr�0-V��	|�Z?�\)\����4c9$~|�h,f¾�b�u��������O������Q�j<_�
��b��!�I�J��F�\ӹ��p��Xĸ8\,�gx��|�&��E������(��#�h[�ЧX3�S��I#�7�)F�%�fI��2����J�p�^�~Yjy�+�v���kK�R�	�&6B�l��'R�]w0�}�k님�.���j�������P��������%{���o����)��u��(�A����|x�J�\f��^F���d�u|X��S���@�O;;�e�����9�������ƆD�c0Q{�b�U$��x��� �EU����b�</ҫ���$�㋵�讂)�̊J]����C�yu�0mY��mfT���ܒ�����*�N��܂٠�;�'��ô���i��������
��7�ym�QF�(ڞ�@5կ�YE�G�m��0���:Z��&K�ӕ��I�_o]�ʹ��mO�g�m��Js*�MqIȇr�}��/��\�/�	,"	ʙ�H����}V�.���Ԛ� �����l�E���R2�Ǹ�99����tu�5�"KR���4�S�� ý�4^��M$��C鑀{��1�����hz���O��į,��4����1���w[�q/�Ո$�5�۴��[��Og���(�OnO�"���/��[r����j�2=)Cx\:��B��@-"�	q;șc�@L��(H�#UpjZi��=Z<E�l�er�
@\_F�>=�O�Yv=���,%X��m��h�ĂE�fNR?�MlJ��)���П'�8ew��{�����Zx �0kAMK�C(� �O4�ۊ�v�{6u���#q�����v��$ט������[�Pmo#Pr�o&끬���t12p�3�I�15��w&< }QK���K�TO��X�y2��w��N��kә#d�U]�Y���(�����$i�kB�5�_al��ܦ�L�����V�V�vx���F6JK�ϭ(Y�,#v%&�Y�͟uOy�G��]���d��"��b0��$���'�gU�i���]Ȭ!�|r*��DTDOl(X���x=��63�)��^m_�ڜ������I$��/Yl�6���0�BǮ�_3D�|،��"�W�pb�˷!���[���[:���A�7�4B�?�챳~� a9I��ED|���>��mF�T��$���<�Dq5�|�57���Ҩ5��K1���ͽQB��Oc�M���T����H��X��H�LUؾ��}���jR�X��C�X�w2��Vs$��"!���݊?^���p'�q�=�R5�7�\-$>�;��#��O�Nz���X�b-���`��J<C��7;e`SUb&��@X�D���y�j3�jEg�ߪY[N��
rI?!�MF�d�_�K+*=Q������rt�&51~�r�}�H�\K1�KA���·ů��yH��h�M�7��gs��5R����� ���d�J�T8N��]���g
z3��E	�_�����>l>l���80�����<]��k\�u~���^�y�&��O��
%���ǉ��� �*�A��#���߹�������}��l�SȾ `��>q~�f��{�F-� *: ��_��Jʚ�7�X��p:&�I(��0�d���x��!�A�E
����X[�����e�<˄8O�%pܪ0y���6GfL�l��9_�!����a�aw^�A���-%�W�`����3��Ow;�RWUEj��~����D�>I�G����S%	U,:"k��1�V�C��S�>��}þ�m��5�-��>q���b�밻��[�)��d�6Ԏ�@H#��W�RUɿ����B�������v����؆v����:���B�y%z��KU��0�����;x!��-<�{��9YY�	��v�-��̘�j�����*+�Z#�Md���|��u���@�O���F��X 	k���9�f���◁����������<_�GqF�Nx ٰ���`��S�G*���3����z����Q����LΦ\)�YB�u�EE@k��S�ď��DZ	D��Pu��tR��K�����h��hI��`c����s���+D��Mߦ^�����:&�?X~�c�[K��"?}7�M�/<��^j�[�Oi:ڌ$���
�� ӟ0�PD)��Q4����Wpm�|��ȏR�R_��;S3�ůT�PZ!��Q�����i��)Qj*�j�}���v���c�O��=Q���B����=MQoM����"k5J��p&���,�������6���Z�Ue`z�,�����%Isn���y̯�4B��Q������C�+��5S�^�g�'�s�N�6��8���rr����2zݦ8��ay��gv<(���h0,�@S=�ˁ��#��ӀB���N����>g��|���Yl�Td�'�ڳҷ5��7�6��e�R�S�wc�8��vt��ra�!��;T�u�$�����Χ������v�ֲ4�3�wE�_y}�������)�D�@�AAQx���[�4�,=?�.��0^�|����7tM�A�F'�h�� $!���*P3����h���O�/�kh��OM��sa���wOx~�K!��m�pQ�L�菺V���U!�;�kAǹ�ߐb���g�#aUVt�8u���8���: ۛն���={ԣ��(�裆_$� �c1W�Q�jr����wǁc��g~�㖦��Q����ۍ��Y�Rl�Z�`ZD�i��?�M���16�Aܵ'�G�Et`�#f:�-�s����~ME�l2cTB�D���;�sk�2�����巨���,�Z��U���Z�֓kmg�E�O���,�E�z����.�$"�F06���ʁ��|�nGu��z9���)��cp���@��j�?F����r��r*�(��D'k��G�5�j_��ig=Nt_m/4�z���_ډI��FWL��ׁ��"W��+�;�����f��I/v��eNղ��������b��!DM+�e�mr?� ̩J9m�x⳰+�g��ݢ2<�k4ֵ�� ��?�Qu�ź3�ƕV�҈m��j�*PbN�TrC9uck=<H�msm�)��C���������l�o~�|���ȸ����QᜇY��
�]�1���K�O+����\%u�V��u���!,�T����� ���)9�^�p�#���%��`���׿�]Z}��(h"l2RR�,1H�tDDD��Ԝx���ga8�:�����rɱ�ʮ�@}�nl��O�/�FekTVߟ'.���-��ʟr��&��yo���k�ˋS��F�YK#����P�t��a�
���i��ɺ��l.\��d���*J��=1������/��aM���ks�DY[���Vx~�]�}_�p~ ;��l�gM�?3�5(��PHRB�ި�=ó�m퐥�%��N/��M[)���U�۴Ƕ�<��dYq�?"m*/��`	�E��ۨZ��;u�wwn3#��#�:@ ����$i7A�{o7I�� ~�^����"�?8~{M�ɦ�A��a��Q0�����}��)��=?/�ή.+Q
�g�sk��v�����"F� ���J'A:vOI��ꖳ�.\A>q[���Ȝ�7��,b���(O<�!��>�.�~�j�X����R��^9J}gz i���ɒ����� ��yd6�Җ�1|Vm�~mɹ����K�����3�u�(��K����@�{w��>
ǸN�rX�Rzws�{�l̩�3�|K�.�X�Lg;���T���tt�奫��U��5��s�C�� )�φ�=��D2^���
?�.�����96ǳ�^<��.�I��F���8T�Z��E�a���޳_ݒ��D�ʲ�f��
�qV
}��e�씗������s&Tׅi����nװP��%�m�9��²����~ٷw�����8���A�w񪋷��&ʱ�%	�dFX��M�R�u�т�k�Zw��:Y�`�R��I����G����q%�7�.��ķ	��
5�"������c�.��No��\=y/_�y|���<�@�A�-�6,\�5���4�ľX�B����C�^l|��t�)?��:"Z�.�gB�]s;���!���Q�	�IY2������8����'�<b]���X1������>F/��j^����� {q��m�7�*�¶������J�l�n���ͻ�Ǩ6����F�(v�O�R�����`�E����!q�ܤ�6��� 1�������_���W:�|m�Qn�<wFU5�e%F0ӣ�SC��gY��h�[4V܉Cb�_�d+#�^%.��j�t��>y��A>��(�B��EL0���f�6Kd�Q��p��_pC�f%�c'u�D��u=�B��7�����V�>��ڽ�d�*�u�.2��XC�2I���m�� �� ��/,f���`����
�O��
u`#�v��2���#�s+��~�q�z$��r�]j3��j�}؂O�~�{>\�������J�W8aN��Kl[zؼ�Ź����k���C�\\(���:��\qm5��S�u����p+_�U;�$�z5t�g^޺���98�V9"��RK�����~��c�c&��Z �7�7(n&jB�'��w�H�O��ghn[~
NA�lޫ}E�����P%&�c�M��1�D�),|�<�P秾x��,���L�E�a#~5�62�f,	�
���ւ�B�S�f�&����a*[���b4V�r
[��J��]M��(] �g�w�% d��]H���F�8�@��q(s�J>*�ـ>�\��͘�Ae.��ݓ�>�x�W0-��1�&5�X�̀��"I����Ց�W�����<�/j��Bh�A��v?�n�`z��ٽ����k�{�������vk�}�
��������1���-7[��O���E8a�� x�;�ù�Я�EcP�q���E��P��7�r�+��OvW}�����=�6	1�T��R �7rF���1�[/�$��qH�|��7.� z�J��4s-/!%���RVSF�3[φL'u����Y�����&�#�5��/D��G.Ҁ�%j߀hW|b��N=�v�+p:��>D7��](p�ܺl"Y�;��@oF�q� ��F�~���� �uL F��xwa�������T����G�5e�.�����j,���Ӕ������6��l�j�9>��7�i�3�i4`GԷQސ���*}����-����ak�U���j���Oܼ/{���-e�kbf~���'�K�����X&1�9=z�9�yn4��!n��,�I֎��܄��܏�������ԏх�ڍ��:��=.��`:���(.�'�!��6�2?M�\䱾�~3��F���`�L�D��t���������8$��T�H1��1���\�?�8��H�	_s�)^�|���E|LL��IE���۶�!�~���37<Mr�v��y1~��h�g�X���v�9�g��p��P;�}*�"Q;��&���ݤr����q��F�/�jvء#�8�l�����;�QR5��W�h{����P�	�%EtG����ׂ�"G'ň��
�#A��9OR�)Y��"���KcFD�5#�d F3�k��/#-b��=�)�f�)ԕ_clT²֍�˨#4z�j�sb!�w�R��!�P0GEL�� ��e���N|�3Jf�:$!�g��K��7��l��2�	u��1� R�î�V,�Ա,m�A���_��
iQ�1Ւ�.��{�5�֒, #M��	�,b���kK�_3�%����VR���+�ߓ�UTe��Þ!��`��YVè�F���%o�Go�%E �����]�8E�Ω��{��m~�o��=�hY���mU6U�����Խ�Z��8V����*�� ���[��و�,\Ւ)���Wp�����b�HG&��2J��&=���B��P	A�Ot��bY�w��M�|+�s��!��-�#���~��{9��3ǳ�����2��ղ6�E�-��r�d����s�֓�������J>k"3]�mș�C��w�f"gB��@Y+�n��� GP�
7�I̛�n��{���د��y�Ϣ;�u*�ry�Qw0(��;�8���h;n3ru�&~��m�7-k�F���k�D+�`���n�F�d�� ٥*�}�m;�9~�n�� �몊�<����R�-<�T%L!/���Z3��)>��MC4cx�.#�I�����v"7��-�w�U���L�kni䉕8\��ٻm�N���~8'��l��LL��O����I��w�_�.͠Ҟ��R(ʆ >��g�n�RI+��[	�A@�������Ӽ�W�VT��b	��ou�B���Χ| �� $�6�!?�2�s����$�~Gj�u�[Q���C���:3�ۘ���V�a�a��i%�<_��[�l
���l//I�ߥ�N=5
�۸��u��@{�լt��yw�H*������I���K{�S��Z֙��v�K��5li���A�����i)�k�J�:G����"P�:_�N�tc���z�O�6�Z�?�)9B�%��6()*�p��Pe�N�[J�?�g
�	�lS>�#>󙾹��B�A�~�;d%�2�u���t�����l����s���E�}���k���17~�	�b�;8VwR����3��
ǔН��S��:!�Y��t_�bP����.�sϘ�a��%�zW8���3$����v.���	�cj�W�O2���@N�^FL��9%�YkRO����Ra���|������W�V\�1���*�rR��Mc�x�CI��$t�DAE�e��ƾ��ԭ:^\���]2O�k�Ϲ��6����x@_�9��$DZ�o�,��>|U�2˼�+��ӡ��웸��G.����O�R'�P_�����r����Ϳ�����N�{�Еu�z߿���6����{��#MB��#�\Z���l	a��(�h��N��M>��Ƃ�eu�p�f���Ǆ���$��'��z��Ϝ\r�v�9]�[�dL��f���#�V�o~-w�2���G���¨�Q �D� 54�dԆk���w�^G z(Z���`��Y[D�}M�e�ٹ�����O͞��H��)�*BoΩ�K����`MI�W�#�A�e����0&�
�gw�C���1����b��b�E���#O_��~q��Lc��5Eo�ә��^LX��u3��s)��RL2�bOJ�s�F������.\��5;Dv�'&�+�U�1���M9tW������ ��U�^Y�v>�3%��Z��9��O�/�C���tsQ��XX���(���B��`]�Oøa�p�:���:D����j�7���O�����M�q�^�bV��׽�|�!()�<���]�$��X��(v�ׁ4����l8���� w���Ws-NC��/�um�og����Y�g�0�ޣ��'LA4Sq��, �FD���
{��6��������eb��J�z�����[��}���i�� ҫ�Y6�Kd޴��K�ܪ&d���Ɵ��.?���,6B/j �)��L ���-[�$�-�&0��b7sL��У�?K���q�.�ۇ�4OD'^ �r� =5[�쨼 �đ����_:�<���T�x�I<x��BguB;�/q��rK����GB{�f\�?~�b�-^��LǴ29�>�ޖC�/�y�j�k|�M�M�#�	�9�!��{�/@����g��Mʠh	�Y8�b�O�I���Ҳ�n�����J�s\_��'̴���)�p�±n���*��x����=����I띄o��f�Քt��^,A;j�������'�'�>L��`k�b��͍Xi����̺�蠠A5,Y�Fz� ��e��6^�H�#D}ϵ����ƥ7udf!�;�����Zb�����	�?�^2CJ^�vWs����l�AR��| :�tY�0.E�e�f6:1��!��ReF]@�c�,�6x�ݭ�E�`�P�)��a�G�E�I���=k�a1���
�N�)����Q�}��^�g5�*h�NU��9� �r%5䓿n��S�/-�����v���D:�p%�r�����D��$i�����&��
8 �����CA��t�+	D҈���5���L��Y6��ta����D��^T��A���X���?�z��yhZʦ�x���6�8��5�Tվ�B�g���`���`'����i$��E�>��nCY�`��A�\�������=O`S���˝;����]A=g"9dQ��<�C1�ٯX���K�#xYE��g�jy�7t5徖=������J�1V/�1� D;v��-﯏�C��5�E�YcWݟ0�9��Fu���d�Ž��ar�j�o4������:�鬛=�	w��x��q��測���8����p��'\ە���˰��#��{�C�Q����5U�1.���X���X�D'@i|:99��������m뻇��=)��l�Ko	��?#�OW�p�
&��Q�
��P�v˫(�H���{�O�?)���[n[�M�>}�Jм8s˟�������K����������/1��S���(4h�u��r�t��Hf>ϔ����y]Rn~t�žk�n�*"����21m�f��"A���b6�Oc�hK��5Ő8A�F�JMշ��6T��3��|�^E#V<d.�7�\33����M	K��!�X��ˬ�
Y�æ�L���$�^K���Io1�ۮb��m��(V>�|��L�������=���M#��Ý�e�F,�^�p?�?֓R��v�z�=���(UQ	�5����*[��$ݺ)`,h�)�BO�J>s2	=m�%���z�Yy��|݊]�D�rhr$M"��}bct|�F�(l���1l�$�����\U��}�A�vW�*io]"\�9v	�Eo6�d
�����4��?2��_�~8C���5!4����{,�� wI�Cִ�o?�V�X/�{���y���q�����5X��7en�dF4(�i	�ץ�]� f�J�teEkh�l��T�$���i�|r�Z`�y�T�$�iI8�H2�_t4e[��&	�ך�n�y{�[��-���tv�`ю	||W�&!i���$#pIn�
7�/9���c�	{��R�Hin�(%b��?Ɖ��>q��tu-�d���p�-�^�Q���̓K�25�uS\���?=�`�3�4W��^�"�Ax��x��-��Vph�߷�����Q^����K��=�(�=�V���IlYG��Y%�YX�
�O��:	E�j�}$
�V�˂R}�Bcjz�^���SJ29�v�ϳ�c?6�}o��yET<ϝ s����4����[��ڹ��L(��\�\}��-Jt[��.L�=5r?Ӎ��}=��@�����?y��Jbu�!�W%9��o0t�ڷ̵���l���[�����~y��+Ig��H��Z���ƹ*5N0��jI�.,K�0�rV�K;�ke������-�s����H��&EJA��T��3D�@�����E'���P�Q�S��4��L��#���%�����|����E}w�rҫ����b�iw��4ߊ�oFe��L�bL��[N����	&������4o�K~7�]��*�y�������).⑄���h�þ:�#
� zA[;1]�݋�����`�[a���rl��'���c�
F��p�$^�k<**q3G��{5�֙AJ#^�D�Y��E~y��q1�'b5�b5�<9$�������osd�m���4u&O/o��1�=*^��+�}x~~�^���]�?b?�vЖ��W�^yI߻4t��Tǜ.�gƾ��!�F�JE}h�|/p���R�����ʏ��g��si�p�V�|�Ʈ��x�J�����"��g���y:�)�f�Ϣ
�H壷�E�]�� ������
 �0?�fǠ˱���1N/�=�Ase�Ϋ�%�W���W+�;Y!��w�RE��\g6/�*^��0��[�����Ds��	{8�vY�Ù�*v�zL ���8^��u�Ȑ��۟����@�W׻,H�/_+p_.����v�,>q�tc���Gዣ#���M���&�ļ�6��[��s�po�+1"�/.M�n�z� ޸|9�R1 L	+	B�x_�3�#<||"�"�'��1 !6�����+�RWL�bMx~*�66d�~w�hb��*�4k�	Ʈq�h�;� k���������@̗/)�v,6��'@��L���]�u�n��By�&���^�OO����Y�����X��!��ExI�N���>k�Qp�1.���f�3���I��Oko}����o�Ktt����z�6�J�Zt{��.Z-���'�O�d�X�U�}hx�0�X�[b8�/ �bvЬ�J/�v� X���$a'D\�^R��,8�_"�5T3[h�?��W.�q4�)8.�J�n6���Nd�=^�R�Vh�RǇ�ϖꜷ^ƶ䞽|A�aF�	I�d�&�Ĳ���18p���E5��B�����w�~��`�^ �?�s�BCCs�N� �)�atd3@������U�I�e~b�5صw\�0̡H��C�J/:���(_-�Q�%A^CJ!I�K����S��.1	k��Ʈ�x���[
0��7B�j��<��ᏈQi~��!IIM��7@'�ji���<�������Z�4�E�>�|�L��[�Y�ǘu��z��bp�E�<I)Mc����"� 1��3
		I��В^��~NT�+a`�c�>������. f-�,��Xh�,���|�Y�v�^�D��9`@	�=JD?���_�W���1��&��Hi�
�
�k�Op]��F�T뿣
5�EH����4>�t��φ�S��W����(��Dc\%r�)��h�w?ܹ���1M��V#�f)+ h%�_=������T ��I```�����)�x�ŵ�O	{W�!�����,?�����[�V�#�|=�w�;�2�'
��̍�Z��5H���H�� J368r^�dQ[-��� �����鿲b�oj��)T� ��*�XKsը�w(Q��8y��`SB�+��N@���q��vX��`�g�錮 ;Jӆ�j��Xc\}�IE� ��$m~�c,hh��� ��@��`PX	 D����V��c\��{���/g�胢��O��
�sČ?O!?������,E�ϋ�y�C(9B>��%}`dDs����ai�\N��}L�����	a����c�>�b p��g�xΰ+#c�y�b"����..��|���<ؖ5�id2fu|m��!�6��^g�b�[�B*J�ZO���Y#4�~1��&2q�+�`S<�g[��z�яB���r�C�~�T�l�ʉ�B�b7��:� B�s�������	�#n|�J���x���y1:�Al�b��g���&��H;�D�������
CD˫2�W�8�J�����0�h�^��}�z��x����u#Ϗ 
��l�]�B̳�U=V	�cO��J�9_WY��P�/�`����J�
����R��e���;��yFP��A�S���D�ճ�TU�[�����F7�8��=��<]uXT����F��Q�^Z�n�{��FiX$E�;�$�AX�s�wW��w����.��9��9�ܙM�~�!��c�!�Kt�x�(��\NV�o?���p��r�'�Y��l񰻣�J�u_�M�lRQr�7	C����d��Q��#��{9o��4���k�S�9������F�B��K�0o��Ð6������1��49-��Cȴ�9G��'%�/�@Ex���pCe�/*�.z���2���)1�j�v��+8��� �Q���a>�q@�@�YƉ0n��s7��R0�Q��t��d������_��IJ0�D��0�`�Lr�������z���.�2���RiG������Wa�H\�!WEZ�������c�=�EZ?�0ς�s\? �_�Jo���H�]RJ��v���]�pYy9>���۟v��c�":��8��ۓ���;Huw��o  8���"~n�zP1;.G2"�rʆ�4�I��W1���@�+`B�Y!�c�o|0��(�\mE���5cl�910���p'/|ӀU�,j�l�w���R|<]�������L�ae<�#F�P��:1�-�$ɶ2���Ʒ0<��"��G�_���&x��V�A��b	ݸU�Z�#�~������=?0p *EXd#0K�X��2�O���s��Miٛv�T�}�T5���1m�<9ۈ�U<�>p�������XU�Ԛ/,��#OL������(��C�>�񺟾:��~��J� �42�1�����TV6�5�|�z��	�<$�����d6=�F��0��$���BEX���:,�KS������?����_��-��}}��|�vI����a�6���!|����ge(��`��+ܦ+Ъ"T���w�w`:�ڛ�v�p9����µ%�:qJ�+j�ӛ��BL���� ރJ�đ���zx���sT{DC��8��E+�Z�D`hEzq�f5���.����) �X/	��{���-��N�|.qy}t�	�5�ZHx�C��a��_���?�ҿF��{�,�P~��è$����B�����I�aBV�=�V��P����{C|W6�iK�l����ơ������a��w�r�p�%U�997�=�tf�_�b�e�m�#�A���#�w���'PF�Rac'��ϊ�@�%?�2���˓܇�ԣ�h�B�X��R���ϳp~6�W�&o���+Am2��񂣚�~�����;J�m�Nl��~�[(adZ~���V?�h�ewa�d�-�dƞC͍Ӗ_���(ϙ��SÝx4� ��������^Ի�o@r����
���zL-�˭�"��3����}����\��s�}^�]��:��o�����/�:ӡn	�˘AY�|kEe��ɱ�^��������mE�N�"�Y�q��K��!7D$Y	���0��MCk9t��u�>���|c��E��#����]�-�&�x�>d�=���&���wH(�t
6+u��iO�)C5R9�H6Ltw�����UJIgIY����mLcͷ��\Q�e�	�,�;Xr0�GJ����h�Hwcw���;;���'s>��[��(�&P��@h!J8C������g��j�~�բ��6�Ym�ve1�lE���D~y���>��6��g��0��6��7,�Q��,@����
�Wb��"�<�3����~^��n�0ʽD�1f/�ɰ�9dw��hݯ��_�(�܊�X�M�[��[,ZD�|���c�X�2}n�`/ALAII	�S�ݢ��V��$pP�1!.�����Nxx-��/Wh~��௄�|�L?<�׼��]�kp�J/>�J����Z��ᓕ`��R��-Rr.�rr�!?J!&�r�J����P�q>�6�������p-��~{�we�d<�婃��(��*��ͳo'Ȇl��d��Mk�@>�9�3 ~x�8j�=}�8�����N"���XB�q�]�� ��{9�q#��sfX�}���"�R��I��$[�Qem�����v9����0t&��[�꟏T��ʾ����<6���z����Qp'���ѺAQ�8�X�jY���-5�em��R�js3N�S��O�NN��iD�?I�"��bm�<�}�a��2���,�*V���Α��U!�0�ԟ}`��R�ۮ��݅�2���0F*�D���6�*>Q;Ê8�1�s�*��Q���ܫ�%^�_L*5Yypj��x�;̕��-F����r�����e�3\�s��Z%K"}�jn3�O��z�x�:���L��h�/>�Z��z���0-!66v�u/���=	�h�.���G0���F�D�ø�=�R�>����چ���K{"_ݵ�*3��1�s��˦0��˙/�fT=�7��~i���"��ۅ1��ǎ�TM�h�3���}�;m�r)t�"0�\e�3�A\'�"[N�s���[ �S\D{�B���o}�D���6l�V?�!�E���ܘ�Nዉ�8z�k�Qn���D^Ɲ_�ǁY�3d�@�� �4i@�����gZ:�~¯��K~1�M,��Z�>��[�s&s���İLb�Cu���mƓ)�)D�9c";�==;C�ñ�J,�����a�E��7�C"}�?t��4� �+΅���Z==��Jy'}���Eqԁ�gƒœ��I�v�ȳ慿�����s%����~N;jcАqϞW�4�ȋ�j9������8�ZN��aͻ&D�=aʕ�L���.@�0� TAm��D�o����0Go��;�I��z�Q���)��!kC��:�j��
�8�L�r|_p�������׵����<��q����R��p��9Ҵ�b��ȤNA%`F�J����%���iqn����\�	#ɓ�1:�>�.D�]w%	����RNAD	3�r�Ԫb�1���!�_V�%3��=�iRw�^w�b�g�/(�A�ֳ0���v2�b���5�O&=�m:����D����HcD������a�}ּ�*w� �A�4�����ȎZ�T�`�P������II��H
v�_�"W�S��W=rO<V�Ը��L�{q�G~��ri�%�l�)�"�,b��~N��
^'�$���.��������#��<X�HJ����%\�"-W��#M8��7N#�!O&�M�ր�#�թu
;�Q~�Ԋ�Њ��+'��DR�u���h�Wq�~�X�o�n1���x:�'�|�,.PB����i1��υ>z�N�y����z������LW/���~�Zp�0��������[�&�kZq��M��x6H.rUG�����RL[�g�-८��H������>��GF�E���E��S"���晑���g+>�Y��6�ղ��lj%���J6р��m4h���[`�V�X��_qhk�\���`61���Վܰ����C��Ȓ	�?��5�x��5��b�:%�}�#H%��V�5�{�7�cH��Gb���7oWK�_���j2��pR?ϰ�'𢣬T0Euo%��������<����M"������2}��:�b?[��E1��ت�9T(��Cr�^o��8�:�]ot9�����A@���tY���(�wj-�;}B���^DU����������:�=��u���  '}�_��	2���<].D��+�Q� �����=;n�8��1�|�bR�^Dr�4���ˇQ˛Qˇa���=�Q93�c�W׋�A��pOգ�y�Yyuޣ�O|�ӹ̩�z�s� �ޔ4��s�#��
�oi�s�(ZB"*4�ԩ���G�qۣ���yA*���dF6��7��bȋ�u�d�^I�I��Lϑ�hJ��kL��^�W�1�n�n�=&9��,�P�V`��q�$3�vJ2�Q�"&Sf(|���k�)��4���r4�o�����:Ar�bK���  7pm9��u���U��_��)8z;!w��q�W�gp��>56OMQ���%���n��hq�8�pG�<��zW]���HM�T?k4�"+����G�����ͩm�PD[��i�4܎���Ta��;�{r�R���}|t��#:q�u�I�������1�R���	c��{��Եx>�z@�!r���R���5V�o>H�4�������f5�]��ZaUL%2_����!��:����'��Vq�8GC�k8)�������RUnr���)��2�F��N�4������?��D�e"����~�8���t6����ZW��*��	�T𜜈��F'Qj�/��-ۚ�#!� ��l���6G����R�a�eAn��=uS���+�H�� �2y6����Z�g�M�d�� K<��/��n3�� 
laNoo��Y�����ul��0tLZ�+B��혏�n�!J4��QI�q��x���=��)�?E`�c�0s�ӹ�UIf��}'vSq?��~�ĝ�WW��.X��ƾ�|�~�$���L�ɲa�t�(j芀O��:�&bǜ���_*���})p,��t�Z�՜z���_C���<�vx�X@�ĉ��'�Sb�kaa����C��čo�Uq[t���+�g>��Y7؉Q��ZJ�˵b+��1׌[�/"@�G~t.�_N���^���E'j�VT�
�pwx�B���E�b�^���͏���y��DJM9���CJ���`;��:�T�x�d�]x��jY6���`��J�1G^���8rO3$`v� ?�7l��3�7A~�!����;�<q���C9+6~qD�9�ڢDcl3�q.���-� 0�c��Y�C����+:��y��G&UXt,���z�#���ɠ�����ubCO�#���6�q���ZF�c�,�Zjua9�V��h������e��t^��(s������ ��n����d�[9��?a�G�ѭ�<V%�w�ί��}3L�V����`JǾ;����OF@�!H�TJ�A���C�Kf�>���x��pX�=��M�$0�1�[N�F8�ѓ��N�w��-�����c�����z�t8Zx+��9-~n`�G�>5�T8G' j��t�-X���	���3:c�IΩ��;.�8l���N��O.�T�p�ϡ���Tt�1W���p�>��s����t�� ����׭wX�����|�o�H��s(�⻊����Q����K|��[q'V��n�$G%�J1��7���U[6��&�σ~L��
O�*tj0�n���P�\��m@� 
���'y���;�Ċ0t��ix��q��}����Y���3���<�k�����e*fG<l�z|.b��R�`Y�ƃ���Ʃ`��l�{f��su�n4��u�����lϊ���{=�dm��դ�� 8������zE�N�_�Q�"F%�q��^ɾ7?��S��c�a�a�P�L�aj�2�H�"剌��|��h���}羣?��!w�b�y����i�I����PT�AA�i�]l������1ee��0M���Gs� W�e���ã���1�~g�R���5�e�8��G����=�P�1������Bk�%@���v�(��4t5tS8W��C{�A�c����K��|�rD�.MD~ ��hS������~Ӣ|-�3��!L��I�ˎL�R�@;���s�Wd-$w2&QUN����S� �����j�ɸ%�{�/�q]n��H�u˶�̠�:&�j�z,���D�/~��.5�g8l^�Q�:jjN��8�G��Y��~cT� �\�hՖk���ۿZ��
v8-T'����R-}u(�;�G��d���3�7�C8�L������cu��x+�e��u�\ő��-�x�+q�;�
<
=�w���ot8X�{~(�I�J��ԩ_E@ә<���M��������tC��e�^Â���~�I_���|��d�,�;β�6�AG�5�b�j�A����Y�є���Vk��cU�p	�d���?(����C<�$r2����ã�]eׄK����-� `9�<364CMCA�L0ܒ���I����Qq�����*N>$v/����J%��f��=��M.���R c3j��ɐ��kڀ��7�]��?�7�xq,�p�B�G��BV6qi��j�$~����%@����r��|A(�iD̀XY���ލ�)l,D�E���H�hr=�_
���p��M�n�ݞ�$�����q4.Q��13D-�7膄1��T7k��*	�~,#�f��z"δ*����.���w�#�=fJX�Z�<�����6��f��E?�_=�����˙�\���[�!ܿ�X��9�q�zI8Y�px��ʉyKK+E7\�	T��Sq�O~�)l.D�U�6Ө��Q5�����El'Sd��wo���-ى敥�5K���{��ZB�q9�.Kn��mΗ�db��&��C�6.U���)SD� �����Z��FG�-����WP߂�6��R�G�Sv���F�(.�G&����[E�3S���0��0��L%�*�
/O7��Y9�US	���4��yl�F����2kx��} 'w�����	^\�ITO�S��$�^nr������{�ـk�O��ē.��*��xu)��`c�{@ǇW�!mjZ%�v�8ŭĚ�h#BsG��K-���k���
  m��:�E����}b�!��u䟠�̇U�4�S�GW���x"&����r=�ߦ.X��w�C����/�����c��e��O�[xm�Q�(�ZNz��r�R��j�<*k���u��O�"k8�Q?.B3/n��Y��[�Ë|R~�3:G�[M���5�*�<��f_�¼v�Cr�����N3��u���=�P���g3rQ�x�T�ʈ�|��� ��*D��6|�d���j!� 0�[pcƠ�)A��|�i�\���i�׸�Ks�3'��{���P���x5i��7��b5D��s,σa�MbD�l�Z�zT��+�/a�o�3��'��S��tָa2��_	S�RX�4��&��)�IE߻�}B�L�Z�e�^�#pł�Z���8�.~������Ս�Ip�SԿq�|�X�[M��������R�����NV9?�C�{8(�&�6�� `����¤��-x����`���6x��щd����ӭ9͝?�D�!����Ų�)�=�Q�P��RY�cD�pyD�5{L�0�G���e�p�$ż�#WR!��b̏�m�Kxp�E`c��A=o*����L���ǈ�����v�x�Qb��?��Z��`�Pg������yo��Y+wE&�O_�uG�;zb��OI�����T��eL�ȓ)C����`���7�JU�U�NH�߫�<G���nU����r��W�<�$W���	�,��X2�M|īm۶%ԃv����܉����`���'��H��MJ����ᦈ_���j%�~uw�.��ƶB��7�Ż-9��%�����'3��{��8��5UJ|x�����cO�!��x=��H|Ч�IbG��j��TF(��Q����Lt�+�bԊhi��e�esū�1�&D�"�kX|���[�>��X�\��F�W��p>�#�/��.1�q�;a�{���Yӫ��ɤ�ݢ���<�8�\}��䧸�R��4|�TJoӖ��d#O��t�H�f�y��l]��
��k���ebf�C wY��7�1�*mH�'3*�K��l[�k�+9�� F�2����K��*�����,n�X޽���fB�N�WaX�=KƎ&��#�v�O��E�mrDˑ��YrDD�y�;�+���2~�\}�V��g�`���%Q�=��)�߈6�N�A�����3 ���[b���v�z�ʇ�$ү�����lL���ݵ���&1`zk�n������4i%E���lf:#�i��k���{#�`"��O��d�CR7"�6���C�>u̇5�>�3�Y��	m-eE�xJ*�%u#��ߗڐM�u>wZUQ|���v�J�w?�L�ӱ��F��SO�e���^�l��ݲ/�=w��z	Y�?�jS���K~�`���Ѭ���*�wAިo~�,#�� $=��}��Q���KA�O<�bع~w^x^{�	T��9��Ű�36CRlJh{��;T?�ʲ~�ܴ��.v�����!�r~0*��ߕ[��
��Ҩ�m
H��`�pW.�w2I�d]'�p�CG4Cno�kJБҌɃ°�d��ę>��K�۝�ȫ�s�j��+IoW�ؕ����S��-�+�&�(�A���5�j�=�;Ҫ���v���es�ʯ�RU1�q.4S��vV
��aM�e�	��K_m8�UF�9�(�i��gQ�TX�5hsl�)���ũ��.@m��f���1n��b{j��r�&���M�QjM�LU�g4ϥ�S�a~���j�J���]>��%�©��ī{��R�|��z�ę���W?8��W/Z�ڊ1�
��|��E���}��i��>5��4�~)��o���Locrr�/��URk7�O����(�Z��Ԝ�b,�/ȕ�}r���f��T;wSl�v3f��]oY�~
w�����0��^$-v����,ō���@[ɠQU��q�)S�����R:lv�\٧t���מ�G�
���<o����ҋ�4�/�R�#Q�ʖ�g�n<_�b9���4�713!�	���+\S���l��5�0���Uu����cI�D~~iI���1�|��o�K�o�j?�gr>lZ6�Lx��$ ��4�lk�0��{�_ &���|u6����>�qOZ1
�7����&)���� �vva[<�_ʾ�UQE?v�'w\�Լ��v$�z
�E��^hu�!�'�.�[����5ݣvs�^+'��ç��W�e�֡���M�jZ)��\:�8�0��z&*J��H!�&�D�L?���L�2?�8y1�4ՑWw��K�ˊ/4��������Xni�h�B��,6�4�΅�B�a��eHgJP��"�~�|���K
�W[�X�Ǳ��}i�w��\�����
���)TO�,��>?��M�ux_���9{/ޟqa�9W��r��T�7�Y�>�W~2K$.Q?��Y�!���x<}:�I���a��>ALU� Fh�=������
� ��=@�l-cԍ�=���0)7���>r��ЩW_M���!s��zG���]�$�8BĘ��4u�4��(�[�9�U��� ib�|��O�����Xw5���]�D�9��Wff��7��	�� �����fu�o�dT�7���V7Iճ۸���X���֚?g�c�w��Zu;�
r�9���Qm�-$ݹ�nD�]�ϵ��+}ɠ�� "�$�,�|�#
[��]��f�Cj ��Ja.���V��6Kp��	n�����2~%@L����c���������:�,�p�Sݘ~��pxhfp����{�k��Q�nq�Al0x�V^�q�Ⱥ�����O����H�x��מ�i��m���w"����s�K��G{��C.�Y���!�5/dN�[������W�~��H��覾�f.��g��t���TOd�L������	\��y0Y�е�A�)��op#���y�}۝�q��?�=ҋ���<|m�\^�*��q���m=�j���QS^l����;�pL!�� {+M��գ	��4'�I���#��b����U��i�mȃ2�K�O��#:��Čvқ��s�����.�wЏUA'`��������K-ߒfx���xV�����p���~��t��wBȠ�������;sm�׷��SFyʩL��DQ��H��?�{:�:�w4<����'O,j�_6�����J���,5]ܟ��Ӹ>��A���n׎�/�ʹT�l�aIha���y��UI�m�R���;u����+lՄ����|�v���uv{۹���a0��[�M�.�~�F)y9N�kT'M���e�>U1$��(����7{u��s��gu籤�^9W����a� �N�Ѣ�A��"Z��I>�[�<;���S��,�ުP�p\c���lZ:`�F9`<�������y��0 �;�rf5�O@�cJ[VD��U{';�w�G��[��#����=hd���lg>I�l���Y
�(��W*����5C�cMO�g\j�!SzO��*�^"�#�aГO��t3����9��K����_��Z�]&`��Kv���1���7��܆b���:��u��\&�~±<�����l��U$�����n˵��Ec�����	�H(��J��܌c�˞�1���7��Igs;e����/�N��H����H������S�m{� �U"In?��nd�@�23���5���4a�{��P`c���[ۑ*����$[-ۮ�u�%��D�>�x�#Iv��K<>ݕ6R2��v'�m6%ܝ�e��C d:��[�3���/���lo�W��(�#����5�b,��ߖ�]V�i*��rt��Y{��غ�r�G��lʉ�4^�h�����������3�hTگL1�ع:�K�UA┋t�ڦ���j�TZu
>h������K0c��*2�;~�W�q-��$����-��4���甩Y��O��E�@J���i,�	 BB.�K�Y6�~n̳�~r��3Ӥ�@�Cr���Z��7Y54wR~�Lh�E�/OZAB��+��-���`�M+,AWCBw�����׊��Vm�ҜX:��D	cL�)e�3�<�^�.���kQ��-���Sێ}%��eh�p^ʯ�ݚ��}8ᅶ?��o�y]���u�q3���� �������E����j�0�L��u�ȁN-`TYNrTHYC�%3|zP	�~��IM�񄡞��
G�W��/�ͤ�D��6�D��+�B@">�tޙ���#��4;�P]�~u���~y���	��E�q�)O��n�;��߭�PX�!��>4�ϗ�Y�P�4/��k��I�!�^��o�bO�B�1�v 7�'��%[U�����7ꔢ����9��C�o�/�'�;�"�8��jU ;�eն�b�����*
mN�<�lTL���5wm� �@~+�^L�D]i� �N�=�H�$2Tt���O��G����,�*7��sTn�}۫`����,&��:�ej{�ݹ$��o�T4��&c-��79x�oq1�mA��Ns6zC��"�Ê�bv�������kM3B�\k��A�ϱ�*�G��&8V:s��3��r�rf �O�.��l"Cy�J��8oM��t���}y6Y�7��+n��D@����z/�{�?�D/�7��_=h����v�iЅ��!u�Wn�]վ��A�
���đ�0a��4"��g�9���jq�����"�٬#�>��]R�o2�<�>�@���m�gn������ŝK?���	Q��UC�������䝷���;%����Pnp��&����(nlF��l�eYhi�-ڵqOTNu�2�R�S��b~�Fb_�M�H�/�6�m��������8W�a�Y
CdoϿ���\�h^x��r�5��3�ը*3�E˛����KR�Qy��u��L0�17վ��
���OW�ko&����?�0ÀT��_T@(��~��7��i:�8._:��`����;}�H�o��)���'�(�gz��LEOڨ��`9�pǵ3/��\����[c�㱊�|_r�.�u,|e1�M%�68ј�[~�!�cS�gj ���:��?�$�O�Z&��v7�b0n���_h���B���U�p���j�m�?4Z�IY5/��R��jIF��ED�Ugϭ�~�[p�̵���@-�.�ӱ�aE�;^��m-A��ᇉǀ7�Cy���~I ��x!�%N9A<J�GR�?�
������]��������Fbc��W6�9n����}��u����|5aH$BIC�1��(S0�U6�יǪ-�V2���g��bf8`|h�����J�����P�g�3C*w� ��7���"�һ.������tD�R�i�'nB�H���Pm��X ޱG�L�C{m7��qE�^q�x����y�{f2}|r/b���?R~�/�9�O1g��AM�/����H�q���4~�BN�v���}]�0{�`vJ�%Ƶ���	fzO�Z��k���j@����
n�y���vu�	��LM�a��g?��KD��e��7*�bI㬠����II�$�L1۷&|��C�%:cx~"���	�#�8a��L��# V�	��4��g=n�6n�fǰ0�߯ܵ��\I�-��B�y�	B־�L����vi%'g){7vB���]��F��O��<FqCD{`4��}��Bͱ���2�l����tF�s��o���ޛtj#��nL&�O�^� M�V|#��� ����@�.�j15,��)L�	�]��\;�+���G�l>��E�Ok���� ����	Y����2�\KR-��[��)k�G�2����w07�,c!5o�����Rʨ�D�������(�f�.�}5l��8gp���c��\`S����*m��x2��my3��������&�h#���6���[y�DB�Y�UQ�A,��0[�7�ׯ�\�Bړ;�&yQ�0^	�x�� (;�<�3T��VS9\z�0�U��p�ҷZ X�u� ��r\��qg�P�g������<TU��h���v�wWI&��cP-�1yź,����a�(�mC�F>�%- (gn]:ea�8ٱ��!�g���Rߪr����ĩ;��p,���v�������D��~���lI�뤰��EN�e]	�y|nfl�yg�Cr�|<��nk���z~��)7���f\�B�]&z�E
^��׌J$3-w]��'e���[�:j�U�:gKZ�NȐ��o��?0����c$Q��#����u�?X�f,�9ǣ�0�����%����㈼+�u�k'�@<�o�TWt'�XP`m��^�}2��ALe���L] 0�)��֚M]qfu:L�'("՜���IE���M|NX��[k�ᘟ9����q�m*���<,AS�?�SrQ壚+�g����k���M�e/v�*l����̀��:0Չ(nRCmS ѺS;�Oe#��Uh�={b��<.��}�G��&�����e����
�e+ϟ��>==�G�\�q�)�Mr��ٷ
���Ϛ1���]#�Z|	��\J�)O�]��*�S�nWC��؂SUݹ޳y{�G.ϲ��?��"�7���u1g��z^'E{P�J�뙽�7�Y磥;m��M^_g/����ߚ���i�B�B�#>Z]e�Jqҫ�w$�q�ZIi"��N�eB�I47���-�;y`	��r��C�ŵ VU�y�F�dJ�����5Y����|�ɼ���>�~52�:�E�7�Rsaj�ɧȪ2 f栖]�Ȟ��qn�=A�-��g��o��D��<���4��_�.�w��3�����D|����ti6Y���C����ŴҰUM̄+�%-�Hh�@<f=�k�2�2�Ae�`H�9�)Ѥ�E���T��ٷ9JX�l4sA$�G��Mkz��V"�y�ö�Xl����GҶ� ��֛��d���d��J�cW����7�@�[�"VkP�,1��u�y����;���Gշ�Z��.K"��J�f6���H�1�ȶ�#��}5�(�"���s<�ޞ�d�O���Mv�~��җ��{�������/���f��`"<���9W�2�7��o��7��X̍�|z0���d�?5]6�#y+|�T`�01Zh�8V�}%�ͳ{�i��	�Hr3�n}T-���Kg�:�wB��(2�Aԃ737�M�*�)�^#]�3 `�Q��`8��=�i�)x����}��^lק���O��	�\����?ߍ^�BA�,����:���֬�V/^H�'mZN�u5<k�&�
��39��G�T23�E]a�i�~s�����$zOjӒ�W4+�/��P���ڃ�Ya��˔�OL�D��{0��$���X�טFͲ�~���܎�p�\^�S���q� �|���jVƆ(ٖwCeXݥyK�*w��z�kcP�?)�zDj�z��`}�ɜ�pk�c�$���f-��a�h�"��H��N�=��|v�ZR,�ܶ�)���dlGJo%���m���/�)S���n2�2���d<%��q���D��EF�����Ǘ���,�B�a���Ǯ�ټ��f2~1�f4gc=Q���s��xd��"�i�=#-��ϫq	����{X`|�^`�-/5��%adE�������ۄ2�i�}�Z�$N�ۘ����x�E_`dSN�������[����;�D�T��ӵ�l�R��P?��=d�eJM9v(ô�W����_}K��T�?Wf�_̬�ޭ���*f�w?Ҳ\&���Ш��Ә��=��L���=���c;��8<MԠ�S�o�ɶ>j��^O���/�ѧ>�L��a�3z�5���!��{����e��a�T�S�0���g˜t΅ɻ��>��6wF?��PJ�	�JR9͡�$�>XI�+<W���T�<ϭB����)�]�oR�)fƓ?�rYQ�0�e���v��/��Q!"�99��7f�]��<(�\�����|�Ni|~�t�`#�`����{|摓����Qe��{�ڮ���a~B��Oi��V6pVc*�Z�,��E��*#i����<��������84�0]/�M�:���^H3�?3�}3�{�c@+�R�b��ݽ�}�jvDeT~�w���>p� ��2��o<���%����m F{�5���`����j+'?[����qC�u�!t�<j���Q��o{��,�/������m�N O�����̈�� �,�2�;+�C���?跎�~;L����,�L�E���PBeo[�v�o�&TI���U^Ni��O�	 �b&��ٴ~��1�M��)aEsz0b(k����]B�9�c�z�,�Wx�D"]�~g�S�5��g�%4�ᚨIbg?\�1 q��ͦ��7$]�Of�<��{�|��<��aEZF���ί8[�'8����: ��"a��Kϒ�/�G8ju.>��8C�r6�:?V�E=�?v�R�����
:V^�E�=�H~}`?�_J�}�g�}'��_�xT@�ctS�<������Q���@V$$R|��)���<����� ��cQ��R捾ʮ��ߙ_{O)*\E�u�.�=)��D3ؑ^��(�r}���(WnC1��..��B�'�r��"DѕF���+UC�C����@s��+��q%^��<���;�֯��|�>01$��n�;�AS�M��Aţ<DT!ӊ[=�7k�$�R���l"ϊ�a��c��Y���D�[CɄ�vJ�i�Q	�m��&��@9&�?h��W7�={���^$LY�i�=�D�zd�{����(߷��9����Gug\e�v=��R�ν���O�0�(��5-r����:C�<�ޏY��ƺ�փ������d=����.�D�O�w_�i����0_�ɚ���4�����܂f@,P�f�!5?L�}�ՓE<t��r�լ�E���z��� �7��:Kr����1a��z��.�|�%joy.��v�h��ML�U�Y��@�7\�����Ję$�n����������A��^+|��B��_��o'�%�l�}�^�(bң
���:*,'U����?�L��:��b�t>.Q*-�S?@O~b8�6���d����u?j1�Jj�V���U�}5���,�����2����{�Jd�ٞ���"����S��դN�AE�v�D����mR���H���>3�[N���Ӭͮ���XZ��ݗ�y�i=1`�!�ظ2&#��%ip3~���C:�q��w$�IwE�1״R�"�8w��`������m��~?[�ܬ�46�nܾ����p�9����V�qu��U�f�W�oÃ�Y����ՙP��9\�X����S�`o���p�.��GU�9�0Ύo��1�O�Z<��1�~"�l@��j�^	pP&>�b��z� H/���e�Á%�fd~��?=S�,�q����s�G4e^Z�b��BX�vc��ֺ���[Yﺶ��/��1����	�](��,1��m,�N���p
����5�;��+��<v�!�)M��8Ȓ1>�oճ۝1�L�h��ak��&�^5���}���-�q�,T>�I"�n?�)�L�,@���ؗ,r����
��
`�#XQ �H�*&��D'J�}�	��B_�����^L�	�RKؿJ)�$��L�!lt�ݬ�^��+R�%�"=1%����m��\/n�X���[кK$l��N��RS>�!B��RдB�{6��]�۟x�U��]��=�k4W��O�7�nS��H���Uz��UDdvw�@��T�Y�*}�cٵ�����Z��coc~��ad��^���w�\nJy]�yfMm���o� ���'��
T��0�]kU����楅i��r2�]�Y��V�J�#��4z�;\�Yj)�;��Y�=(��^�c1�JOt�2]P#L��=�ظ���:���6��6BH�Q9%��������u����,�p[�<ٝ&�Zr3s��U�m���D�������q���nvM��* l��cͲ(���h����1�;���
��mtz�to���#��u����Z�ޑ�N�>k�*��	����lX�}�W�]�ceC��1wK��UD΢f��=�ܖ(Dg(ߕ���wR�eۚ۳�FX�+�#�J��v�
4#?(����B�i������խ���nd1K��
�n��������7�ի����㘉�Wqչ��Aϳ�_�|%��+�Z���W��Y2�.�go�5\�p�w��7WG�R�99�-;e� /n������Q�{�P1�ը90*'��w����?���-����ni$�KJ@�AB:��a�ni�eH������!�j�����}�;�3�:���k���9"�3�m�:&�wxxͻ]����s�b�xBX�pF�k�"|�b��}�|�g�>�%�΂=�E�'�S��n�ٔ�����]�O��ĳ�HlTPG��w��VP�l@��@��t����tz�	����_�7h�����6��+��Nb�dak�ǝx�&K�v_xJ��:J�.2p,$Ҳ�p�����X_4
|f�1-��������o����C�Ә7�v�;cK�;>�rң���Q	r���@��J��2��n?!P'��*�C7�A0�#%$�A aTY�����VQq�Ft)N,C7�ǲ������%��� ����\-��B�I/�����[CL)C	��y;Ѕ��X.��(�5� �����"�u�AA��v��R�v�A|[T;ٳ�M+{�g�uʒfb��A�vZ\��������X*�7��,2m{��Fr�U�{�Or�0�y0:���Ȟ�S�n+���츎;�����2c�U1&(�*3@�8�G�}�6�^py�f�]u��q��zaOY��h��F���Ʀ�{2�����#l�m�U@�>h?W���@7�À",��y\�g7#�_�ĺ��lB��Ck-¡�OI�k���\�{s�J)�Y5~_�{#)u�Q�\�I�_��G��'��%c���+@ڤ,F��'����*����3��w+�y
��?�"�x��.�{�`җ�}�1Ok���r���װw^�!:�����+��67Y-'UԠ�mz/��p۴�hr�;E�S�v�iz��6����.c�b����cU�~�ɳ��a�M���|��c�ɾz�P9�\P�E/b&�΋Q�V��{�cmF'� ��wy����ۂ��0y
W�m ��M�g����?{�����Gٶ�6 ?�}��eL�z�B�kU&�R��^:�+�d��[x�[8����3����ُ��xx܋g��0Y�yF%��T�0�T��/��Y\������p�F��elv�k*&ç3���'	ϡMBoŗ���z���;ڿ�0^�����NI:�
���5�el�9(o���EgM��F������ݑ�s!k��o�;{�?
ڀ�"��:�ñ�������P�X(GG�
H��}Ds�4�͠M-�F�ҴaD57v^��A��8���� ��L)a��S�H@�����s�㫫(��deޓ_�`)}�7�`�mv>���!ΕU�1����<��7ܳᤶ�B�q�� �)g����"QR-�JE��5��n�R�Ú��������NW3��Á4�����V�^�x�^���lȊ!rxK�<[����%��܉�Ă�������3�F"����k�?�~�q)jZV�P�౩�ݬ�_y)iƆ<.#!�ƀ�_H�����I�_d�
)?9#���������sj4.��t4?�(ͥQ�B��YM� ��i��>Au��h�|wȩ΂J��ɕ�ٿOF��,.t�����盾Rف7o�'8�0��JPD�y���Ap������J|댡T2��:o�m�HSߠ%��}@�Y�l���/����ا������k���i�:Un�9!��ˡ���.�9H���ż�b�o�|}��n�,l�un�)��Mt�8YOU�쀂��!�R�V9��7�w�E
ϔcK�Z��a�Ǘ�e�Z�Z��!�ڧ�t?V��ȫއC��ȅ��{E�z���뺈�wh*Zj�v�����0�OL�8{��oY7u=���^�'�G��xՇ���7��;�6��d(d=��������̃�8�|P�Q��^�f�)���HWs>߫��r>Ҹ�m����qBpCaG�Y�����"׸��r���n|�l��#��,6���^�z�]��5Y��K����es��)��	|U��D�����g��}9s���v��
�q�_Aү��Hb8��A�hE�2o:�� q��6�T/��n��*�9q��������7"�D^F��\N�.�/��%��k������7E�*�H�Op���fR�/@↥���"��fm.}��=�����C�Մ�k�A�M���V�v��sq�iV��}�V���[�+��"S��M�K���-�s9����p����'T~�&��C�s�ED����������W����%$Z^rʋ�wmk�A�q����}�*M!C������޹���Yd��++��Վ'p}����E�H�P)]�;E)w�	f��¶�*r V�_�Y�ev�8)��V�ㅯ�e��F���֕BG�JS��g��!y�q{���_	���xp�!nbmͺ�I��A�G����2*͘C,?M�7t[�Q�_Y��g���#�����\�z�"3�U�7��K�~ЖZ#`�Y�g�i�׳��^~ݦ%��:�=�6�EK��8ѻ�uDM#��F�&���K+�k���!�5m^W�j%�9q�������U5�f�L�0q��#��-������MS~ X��� S�t<)!=Ug8�!<�����4���HK�׺zO��0��Cl3PA[L2Y���VZC����C�c�xp:���-m��Ug�x
0�5�F�-H@ƃ7+��\!��6=�hm/�9��h�ϊb�u�K"G�8M�����2'L�T}�.��A;6�.n�a��,(O������X�H_�������p$�� mB�`Aw�Xg��m�Ut�go�x�>;ȗ{U�ז0�ô˰��-L��#y�˒7�C�)�`�`���F.)��y#m�{���� [c!q��\7 �)�Њ��`+]�N\����p"�����j�/���88��\])���2��Q���t�`�ko�`�i#O|�"��4����D�ۄMKrT��j�Q���K]?�%�RH���I����K�n�5l�h:��|C5�}	�l.���Ÿ��=���O��,8��AH�;������ma���5��<��	̋3X��(Ն �c��p�p�M�����ݗl��z��o��A���뾷�dX�����d�T�A����h��^�GOSx�4j���ށ8�CK��W^,��L���ǵ�7���!��w}��KP�L�Yӈ�7�ڑq[!FaqYd?�3[�v���t�Wɑ�$F}��:*֪;�?qB����]�ټG�fW�����Pe�jW���������k�N��,O�𶆠}%y�!�AR(��3�k7�%��ȑ��_�.��t$#�%H6�g7&��8(����ߧ��1�멯bwJ��X玨���cP�o�d�=Û=�CEӅV�Uv�䛹N?��K�C��<��b�y[�Y�5#�7 s4�g��{B�������P����z�V"�����Ҝƻg�ͫ1�=�����~t����XY�����t\�xGrR~�y�����c�ҷG#@/���^X�����`���[����+ʙ8���C��C+��E"\�8঳v�>'h���A��b�/��G,��E��Ň����X�I��.bǳM#�ܪYk�r1�u��u\���~d����K�m7��r�K=pQ(�Eu����rU%�D^d\�2�0[�:T������3�:C�&�d{���k@�j�S[ �'l�L�XQ�{w*滅�8ޠ��<�!�0��K�Mp�h`�4E<˒孨C����Zw������]��L'�k`�C�a��^t��ɀ%�1I���A�#VՌZ6�8�f����J����;��cj�Y�K��˿�/���Yw?��@$����SM8�6x_1e8����������/�(��Fֳ��m���}�">6�t�<�����II�]��,�*�*M�
�i�<EHu����{
�QNb��l�5|�{x�h����Q�0gK���®�c~G��8�VO�3Fo��}�6��ܯL�ނ��n��J��z�ʐ�Y��\�$H>����8�T�|I�Dfg̷?����eA�" ���\)O��C�,�c��e�ʸ!$���:Դa28/̍E����Y~J8��3"x��X���g֭�,I���-�ۓU>��t�7�b�K�|J�K=��J0Y Sk��n����D5����1ōk���7�A�u��S�����~��Tm�&��#��k�I(fՂ� keш�c �w K�w�Y)���p����2�9�:޹�!�v&6�*�=l)���8�v"&z(��ަ�Rҹ��,��Z��zx��ћ f�K�M[ַ�R����W�R��h����w��9�_O��H��!��c�1�ȄV'Y�i=O�µp�u��Ԩ�������;� O͠`��}0�Cf�VF m�������R�b�S�6^A����ǫIn#�?���dK�F���,kK��|5fY܌�������-�6�R�0/��]Z�	���RBu�� %�S�>��n鍉׏Żq���@<�L�r�0�y�g-���QUY���j�ԡ:z�s��A$7u�sx���q���-��ijl��,6�Mu�7��f6��֐͠ӏ��$ 1��R"�m�!�Գ��<oդ����\4����픍m�?uK�/�7-,'Aw�G���-���_��Xs� �<�C��U���D�2�Z�s膴}�e��l#yѷA�W%��&�ڪ��f�To�gT�Ȟ�F'���-"MH{lc�UΨu�C��)��H������� ^V�&�`MWQ8��Et�;����N����"[}|��ul���̴c���x�4zK��y�#�)����z|P� �v�v���9��}%<�2��r������D�����ǧ���j~����M�=f�\�+�'.&�[���ׅ�,�5�<N;�1wR�όA�����ϟ}���luKn��x�~�Z܋=b c���P�/��
xP齙Ș<����|7v���L��+k����)��ó��~	��Y�E�Ց\�8��@�%���i��X�ú\����K��jJ�*S Q̇�B��J�����*t�c��ə�|�aNA��>�ǱN�m)�����!��8�
��b��݊%���k�l���#���H��� �fT�	S��^-�Dp���e2v���n
 �(&t�Y�#4%FLtP��#<�dȚKQ�9\w���u���X���G�Z����|
��u����w1���m���@�ݪ��;��@[g;�Hj1�3�b��#i����1���,�`,,|�E4���wO�d��j�#��=}x�a�k��.�)5��<�W6����J�}ZJl������Hb 7j5zoդ�>�L�����FG[c	�yA<p{�t�H����J˓�_�͇��F%H1�ip���ɃS��ꂊ�"������t-���R�Ԅԫ�5Z��s�c
<��Fz�I�~���K����%�Lkk�}�����������Y-�f��ޣÝX8	"��~Y˴]�~��S��u����i~����t����KoFP��(n�+��շn�jD7Z8�oi����hn��BR~NA�t\9\�n�^��W\����E��Li���)�XԮ��^�ԍMH����Xa���b{n�s�3I���H�S	Iű@��f:��@���`�%7hv3֢�)o��qv�E���RF�9`%�Y�M1��7@;ܚԐ���Ur;����D%$���dH�J�F�d-~��>�!�u��P%k��#C���Nx�)���[Z�M��v��Y|,~=��SU��g���#�Th���6���f����U6e���m;@�`v��Y�̻^�X�n��y~�];&�˲��bAt�z�^*��Z'��`]��>u^�9x���\�r'P�����1�,� ·�wZg� ��&�Ê�|&�Ȓs���3���Y��2�x�w����u�	��j1�_C����tw����㦕!)�%¿6�F>��u�NIȐ$U���"�-/ף���
v#���K?=E�D��!+��q��c6y�p��;
 �Dy6@�7#�}���#���.#��:ݼ���Pe;y�4����$1v��/�����Y�`㩹(>>H1��	����q�;�	�?�ZdT�긯��]�������X�����$�j��Q	rg�@F�ݏ�z6��nRW��vLW��J���.��U'�E?��λR\Vn1��(Ũ3VB\�,�������W���Tk�������zu���Z�\\%�����R���.*��M�cV��!w���z)Y��ض���@�W2��󕕑���jj�o���1�R��&?|v�VN�>�LR=�Px)ZC��w�o��"Cu��}!.�|D�.��iv)E���P�C�8���H�a�l��Þ�A*:!����B�+�1�ky�]D� ���q���T�Nu��52���L���Y�E�!\ #==���/�C��) ��^4���V�����72�D�_??��
36��KÖ��לl��{`�)�yFfO�^�~������C"P��3�7���Z�hV$��R�;���fR�KK�3f2����;+̷#p�LEk��O�F��(�vs���0/�Z�����s���c��"+�;?����R����.as��jQ�M�[�nu�ؘ��>��Y��1檡?�����J��wd��O{�x��)�;;Ч��m��v�a�۴p'"�<�Zu����{aD��c�f28�����Ph��;'�̑׭�^CE�T���(ڿ���I%6�+yS��ܫ.u$�k~�sC!+����*����=��9��k�ꀚț]�G���yTX���o����J����6����	�JvFP�y�d�evz��D��a�O�S�D}my>[��ػ��\>�����o�8&e�����1JCW#$��m��@f�g�C�j�E��~��Ȋl��n4�Jqέ�ʨ�ɖɏ�sv��W��(N���~�۲ ��6vU��U P�*��O�ݎ�n��W�M��;fU�4�򥴛�kSM� ;,�H$��A�Ϧ��:z��c�e�5#���n;��i�0�=U�TM����u�s>WQ�R�jDI��*���`��i;�w[}�(pc�A��0jǅWuN�=�o��S+�I��͕��pn5�����,�w�e�82��>�AD%�$���n�9ѯ��w��� W0�X�-J�r���E�ًofe�7�Dv�[i��T��PX%��f�^]轛9D���Q�kb3��}�B5�߸�zV�m'<�҈�ߐ�ԟ���P$�\xt���2�J��!�,�#~CA}S�<\�����7{QC��&��5Nl�2�&z/��d�c���>�I�]�Iz]��(#7T ��e��[/*����#�oD���c��Jؗ,,/��|��8�+(37�%�%�Ԥ��Ÿѡ6a�v�eb�,*|pu�H�t�����᢬����K��j�(;ٸ�&-���NH�$�5S��+Q���������-��e@����J��VP�f��H$FBU���_�����{��3r���A�����KMw�֋�� ^ݧkU�-0vKeKH�l�Š�|x��sJ����ٶvbF&-�����4�e���N��1F���j���W��s_��a	T�p'@o�x@F�#uӞa���(h�jʺ�ax߹H��KRS0#A�7�Q�3��MS��_.��VD	H'���@]���\�ϴ ]U%z�ŵ�1�{f#U�A;9O�"��V�=b�g��K�c.��H{��?�!Qgg������x�ޮ�"�L�����MRh�K�_"he(DL���@����x0�..<���a�!� �`#CB�v@�o}�:?�xT���J�t�5�9<޲�U8��[�?u�R���|�Z��#��r�උK_z��(f��c��eSKo��֌�Β��h�y�,�����W/� !��(�2�������5�^<0�<8x:�L�_^m��f1-e��@�:���=���M�����nˑ�X�"lq1�Q�����4����ھ���Y��1G�LRM�f�#�ί���/��"��b����JV1!�7�YO!g� C�$�!҄w�u��(�2���1���D�:��/��I��d���d��������G�YR�����!�&R��:��G� �p�Z�}������tl)��#��]���{���H�E��?G��=E��|3?��2@��>*7��������v񬚯��Zu�O�������~FN�ne�!h�϶y� v�Gg%���l)Y�SK�U��mPO l��:'�����)���-��!RT�]O�o'�yw��f�/�Y��"��w��aP�{�*��r7�\��Hb��W���O����Ѻ���mx�+��R�A�e�@@%�6&��+#�0����a&���+?�]�����y=>b�]�f��\!�v>���V�E��Ky;c���9��[;A�7��j�i�X����(����\'��@�Q,�x��[�}���m�zx}	������|��7����X�l[~H��(�\5}�A������ڜ��h2;�rE��`��7�.���c�9���~�7�&�;���ᒀ�
�ɣ9.2�<�X8����o��%��_c�X��W A<���ԗ!{�ݍk�����C/��{��{� 8�{S_a{��}�u3�Y����x���!s��u�.P`_I�})����B�!?��'�n�ZK�m󉔌!�_A�>�cT2à}�O�b�݅�]ٳ�8�:k���G���S���+V��-!�w�j>�KYz��~�D_UEF�9�=�Ũ\Ԍ�'	��|a{]:�*B���.�J����-�74:�I  �W��س\O�D�5����b�r1��CUX�
v9p������re�&ޯ\���[�e�Y�*��[��P���q..?�����Lp� �Z�$�]rO����Ux˦k��'�!��rf}s�M$�§��K���v�Bq]-iGw�UG\0<x�����'��b�>I�"ށ��pُ������%()�����y�8a̯ 	�o��q�=Q�%��W��d�ϼ0�Pm�X���iw�=o������7}A�׭e�tf<��x�ly�-y遳t���Ǟ���8fh���`is�'�d0I��O���n�:���md�+��!|�u�eJm�Q�^�~(�YBoz�%y��Ǆ2�R�S �Ht%;��'[ŭ����u��'W����������-���b� ���,K��F���B�ꍠ�$F�U�����]�l�DԶc&x��S�C~�cB���	Dj�@yR~����G����62�Һ%Hƙ	U�-E,.u^�˓q�)��-�0+��3B�/'��t���vbDN^��DK
B��_���Kv�~h��RAb)� Ec��U����˂fRT��jZT�BI B0��QS�gN������!��9��@c��\ϓ�%��[}'��^pW�LKJW��l�����R6$�޹�bG���eՠ��d�_i��Ŵ��6e�$����6�0�l��������ݴ���b�B����9S��J�]��*�Y�i@!����IC�$$�J���\Q��0Ќn��g����Y,�~7�@'���W��hDY�"'�(N�OB�E=a�b"�~��N3ޠ������^T~��mh�)��0�h�i�M{�����ƨ��s�͚�߳�LtK륕4Lu>5���|-�f��wa,_VP���m�bBS�������Ks��������iJQu��J&��g���������!��V�z��!5@�>�M?�8=�#�w���*��ʳȪ��+�^G�`R3U���A��͗�Mߓ¾�2=��x��w�"�ZXG��l���v�+6�
w
���߫�h�<�����������^�B:]���G@%�ձy��#ظ�lN�例�b��j9�#E�EH@�̉�aݠ⾆?k��-����(���\�a�׎�d3&h��~8_�I�Z%=�З:H�u�%��w93�)�I��5���&H�x���?�!�~�Z���Lƣ,ĺ���������M�%x�]��"����W�1 5u�c��w�N��O[�;%*J{Js�Kqr��*g�I��8�0c��13��0|["*FG~��s
>�^�T�ElE����f�A��O~�A�Ǐd�i4��*5�e��*]�Y],z�6�?��+��{�	k�;�U�[L�$/B�_�۽�����IH��z*֠B��$�?N��ښ�F��<�@^C��G���8Q��L���͚n5�J�/�V�
������}�vǖ�2��!P��Ƒ������'��2;�!L�u�y��^ko��렄	��5�/Eb������q4���0���J�=�ѥ�< Au�WJ*a}!���v���QR?���:4��ob;�����X���)�􍼁r���!�����+v�CT�ú:�'�9�D��j��z�#��	8�7�J#=�IY�0D�/ߣ��e���liû>���ikr����J��}?�����ڒ#�~q�V����=��~�S�'���/��$�����Fe��-`;�Un��,��(��|���6=�U���-�>�#���P��&���d-�C�� ݿA`����s۲�󄁂A�u
�����FQN��5��Df��n�^�j�}�Kk,�Z�d`���p}��S�����Hl�`�x�~��N�a��u]9��5T�<��m����y��(�H6������_�����*��[zށO0h��W�ޡ ��-����Y4�s��+
���_��`��V���<3�����1�%���1��#���n�	��)7LzHJ��F�z>x�.غ&�e��O���]_�NM��r���u�&�"!sQ/Ⱥl�Vn�~/O��	c��~d,�aq��y�V~1p`��K���JH&�lqѵ$߳V	����48T"�ѥ:o��(�=���]����lj�_��V�G:=~sx�폹WatM��]��p(Av+�L~�����L/B53�5�������Y��b)ј�����K8�`����;PIPF��c��70�k��i���f$�hQQ��|�k��y�#��Z�be�@Ӈ� Y$�����l�P�����ڑ_�5� �1�S��"_�������R^AJ%;�Y���%WPP�@���%�)�'F-��a��6���q������'���2��*���,B+C7�iɱ�^��е�%W����P�,������%.���k�y,�G���w�k���������\V%���SM��M���癥n꯸��E0� n;B��RD��.xl�N���I��55 �-�����	N��Xk�����@ы��W�s"�_�|FF�8��x�Tf�"���:�>x9��p�44��tw����J���8�I��6�f2�t�6�*[>��E���yɞc�i|\�r�R���!M���2�jVzr6�D �ЂxX$�(;�Ó[v-��@�?�]��D���ʑ���KB	���1�˥;
=��<0� 9�`�������B����)�V�߁������[�6���L��#���	�kS����hƠ �н��]�;��g�oZZ��c^�y���s��|���Mȕ�C�'�]lYC�:�f��9��Z�a��جu_�
�i��@���N�>��K�޸��\��2-�*�����u��lpO�ݤ�P!�Y�C}�6.Y�-��^�Q�P���D���-�i,��P:8. �6��t��3[a@7"
�"��v�=�b<���LYwn~� S)Jm-���=�az)UJE�&��Fo�3�QR��[*7�æGK~*h@�ә��J��r��=2�b�:gȌ%�l�e[쯭3P":T����+e��j'w�y*<>�G�'<�Hb� �4B��}�`����ڦ�ދ���"Z.+��r�S�ڮ��W�g�-�����@�C�]	<��X���w~�닡Y��<������ݐs�Y���+���kC�Ƌ��Ձ��e��l��C���{�}�4J%G&���`���'�[����U���s�9�,T\�cl7@uųQ�թ8D"�m;\V_�I������^�@��+30�eB��jR�5�W]�3��?�t)���=��/oЍ��V~#�!?>�~����E�^��&� pg�������Qo��T�����;5[v��Z�y`2tfV�����m��4��m�$V�b���Lթ�#rWQ�������ѻ�b��êԁk��-%{���L��L׀�C�62�B���s�� ;.d���+�v%-��5��&�S��
r��{����;c�;���f���>�<�P�dn{�즟���U[����C2�'W窓(R�B4�棟�N#�1�0���6X��B����2��s�N�a�c�N~HT�z�/�%�A_p>�6�&��z�4>"�ϖsL}7���l�GJ�c��6.�R�K�
������UKUO�*6�gg�&߾���4�S$�][v�wj9Ns���y�Ѵ*�.��eWXg�(�r�u���w����٪�^�(��8�Ts�Z�hrL�]�K�3!u���wƧ�e���&=��S@�>�^�?�
�С3ҊW�M5C�A��Kdױ-ױ=����E:q�ՅP��Cș'̺%�����t����ǭɏ�^k�m@�;W�&����h8zIV����DI���/�w:1�k�A�=�;y}� �m�����m���ah��0�e����j����Z�-��*�+�G�(#��T�]��}G@�ܩn���@�b��r¦��:3\�=&�9�6�ᩋ(���X\u��Gc��r,��|���@pm�Ӌ���̈́�_d����U�m.�wO���#5.�E�;7�ރv!w�N�����?٘ ~���ĉ�g�:Ȉ,Z<{<<U�����~+�z�ph4b���`W,���Q��sc6�����R�+�yy�i̇�a��D���E}wM���r��mU���һ=��-�4
���Y���ƾˁʶ�Z�̗��&T��R+�+��Db���7��Q�p��͵卦'Ưt-�kf�	L|j���G�ڵ/�=�7<�af5�,=+d�a0	���OL����b��?�[K� ��	�|�ՈXK�/� I���ܡ�$�KD�D����[����+'�ѳ�zC]ȡ{�[\�t��v�
��4�s���r����}Xe��Z����;���?��3�cS����fc�Z6��$[9x�J=a���j����}��^�_>v�3��2���F/�a����߃�;':_��]�d�M�����sxmGVz~/xŋ��$x��Ht�x�@��$SM] ϱ	_#g]���-�݄x�]��3�c��9O~��C��t�RS�.���c �~g��i�GdQsdzM�_����ŗ�(����	��;\.z�3'�Z*��j.��cf!no?Cg �^=����*d��?Fg6϶��7��?ƌ�\f��p~�ҝ�=>z��|B0�8���k�E��
��W�����duV0 5�����Y�㦍<yt�I�ؠ�ƯƂ��Ѝ���<�L���׽�Q�/���� ����J�ĝ��5�]s�\���g���@��d��9���<!� x<�����9?o��D��O��S`��"����n=uE4*z���"����
�;Q��Գ�)�c�/������6�D�ok��ݡ�:ſ�o"Έ��_���I��=m���?pDG�.�@Y)�ȋ�Qw�<Ί~�]/�*�x��~��;���$Ezq���T�3t�}v�Z�Œ�p���rʌz�2}m����<��ao`�=[���A��M���}n�����$#��X
��(Fz����9$o�T&�qz���<�2������q��W� ���ى���uk�X�����/�LE������3GE���k	-�]`u����js���8}����c���rv~Ta�9AAsZ��3;3�ch�	�G@��o��(��=e���W"�%��z����N&�Fғ��?+�BW��^|�zQtoؠ
H�8��@L��t�:���>ʌ3 e���y}�\��Y�AH�uQ�_�a~.jqR?�J/����Z�gt��������������*�}������$��~*��_����(�f��rt�m�f;eN��ּ�|($Y�e����:���+���ڗ:����Z
z-������nr���������v��+�]��׃��Ҧ{� ���8� e��L�X��g(����&3 d��((d�wn�G������ފcΘ51�pV�Z�gM�~!�%%���X����# !H����(nX6�g_�=�rѣ��ɫ|g9�<l<!�0c��t�L����d'!��J��Dz�#�R-@R���H�ˉ���	�5���g,N�c������y�d��5=z��E����J&���p�ht���6.�����P�>V���p����A�:Z�+@�p�ߨ����Z��x�L]t��>a����^�R3e����K��nX<۾�%t?����$<[�\��l�ܸ���9���N�]1�s��/�vR�lJ��hR䇟y5(Z{��k��(���[�~.0����1&���(��Ђ2%nf<��(=��	�����Rs����s%Z�ʟ�y��v�bfS�i#I\��������%)��e!u�u��:�0q�&g�Uț󼲁��hÈ�6��b��љ��d���Z��[�L�B ��J�����nD��]Sik�TQ��u;*�^�T�9�'���4�1����X�*mz
���]��� �E�/�}�xeL]>z/�+��~'�2�g3<�9�	��X�����,���xݰ>ܩ-b�������iVy2#�|�L�	�r>ix^�y]Ď'+������e�b�w��yUb�-`��(<[G�V�~a���J-̛ݡ?�h4�2���aK'=��������z�<BZD&^9ԆҒ�,���^�5V2bLG��U��`+�lV��,���M��%?n+��l5��^z�5�`&C;_���|V�Zo	�^9+�
']��&~^{ c��CdY��;�m���9_;�6߸���v��ůE��UJa"��c�Ƌ]���y:߆R����G������]�2��׋�1'�S��ve5�ג�%���$���Z�l����wt:'��wӷ�U^LY�2�1�����%c�o~�����KTJ�@H��\�����+S{�S�q��n(8D˅��=�m����;8~ŋo�k���3��ٿ��Z������,�W4:	\���l�+�,d��xw5?�iN��L�uP�v�׽H8��dS��q�Ha�(_�1Y�`/V�c��ٷ�dཛྷ����-U���]X�Z^c�&�$�D���g���N��;�k2;�g�C�v����1t�O)i'�H䳹������.'�k߳d�oS}�P���h�������߸�	w�i��.��훢�:��������Og����:F/�b��3����;�nY_	�W�O��k�����P_ j�r��a��^(#R���۽*�l]���{�ʋ9XԆE{=�U�1��g�MX6a�v$C
���j� ��..�[�?m��Syz.�`��<�����v�ı��_�4��7YVk��a:.^����Q5�:�`$D��z����"VƊ�x�@����H��u7,Ғ|!Y��H4��4u<m��>+�qr�_���GÛ��9�M��R��_w;3!u6��qt��y��1����l�	�;�����oTs� }��g�ҥ�\m'NN��3�}{W%.�b��T��}y�ۆtW˅uA�F�+@ők�yƄh&��_}�i�-�&\�Ŗ�ᩚ7J�9��a+_�_�A�~H�+_���){~e�Ud�@���sh��G��c�Z��7�4���͝m[���-&M>����+���!��G	Q���8����P������W�٠�M�V�u�{Y<��x�f(��Ri�p���&HF�*BN��mY�dϠ2����LWJo#��/(}�7Y%e|��>�޵U�A�˱�C`W��8Jb�妕]MվR�{���b�j�Y ��Uu��.
oڻ~l�wf讶�$H�qR���_�t��U:K�,2I�^2��5%#zݛ_�w��;���� 1u����ק���!��a��g�[����x�g�o���S�l�	�1�>�YW'���yEt/zb��$���V��X
���ūe���q�f�)�󐓭�2g�S����;fW3����~;���ӥ�j�����8T��eW�>K89�h�,,�]^�~z^Vhc�Ӥ���j���~���0O�&[\�z�w0䦑w�E�t��"^�丆�oEd��Ju3!g+��.��qT���n���<��8�$���M���]�q=/���y�נ�� /�7VVΜ�3\S�¿�p@͝�	��X�Y*���H^q�9���۪�k�g�i����2�"�f�Yk+���]0V��tq�;~�����:��5��� a�;���	�J-W�N�Rz�v��1%-��ˬg�W��m�8��H1���{)(@[�)��'�C����k�"[��+�ϓ��p�;R���M����9/���J�/�J�b��a��YDN��}�p����>�}�$�/��Z0�������P5�p˞�z�?�x:�y�>5���%��h��q�+˛ �"ͧ�����W�7����Q�@�\©�r��/Wy��~8��+Wxwq2:�(�-G��G{~�`Ѧ������at{�,j�W_ξ\s�e���Դߚq�k@�+��m��VYm�������V��>=7�.���FD�杋"�x�d�z��q�
�ix�~�?���J��nm�:���>>
�xD%��~�CsZ�,������ߺׇ�_��k��}�hS.��=��?�/(b�j��j�����oQ}_�0~DAR�CBRB�[��Qi�N�.	���fTD�K�[ax����#���\�̜��ޫ��{�6�v.=z�s[	Pnx��fّ��eԓ+O�z��|y�����Vn��,b�<68�	���Ӗ�y�,��N��$9�/2���^h�)lyMA��!�YZ^��4{���o��x!e_kj2�B$��\��@�,q��W�}F�T4�4
0����@:���
���̽�;H�6y	��C1�����[�,���V��v���e�N8�	�$�~r�k�a�t.ޣ�.D�o�'ٯ�k�E[}]�lLIKWx!���7��,�m�g��6�q���eKNJ@�ڶT����-e)��_�a9�ec��>�_�g9����ǭ��#��u"�b3j���Z�wy��]ӊ�!�R�P�����;H���&�Cټ��D���V�Ǐ�ҙ�߄,�Cr����֜�� � 	���(���v��ʈ�����x�@γP�{}�K���%��up�U���1u�~E��~]yEq>&b���7�X��	T�1��s����z�W �6D�ܻ�&�ڞNPT��� �&/}n����h��dI8�lj���R�����Qo�7�cJ?�}I(�Z���<RG�6���,��}|Q}~��6td�p�+ްa���O�Z,��?��vpKE��m1A4ً�?D��u���o&�x�u�oW�Z��d�y���NC't����O��{y�놀�7�	��|��Q��{
Wz��(y��>l�h���4�C�	W��%��W�ټ:���6(�
�R���.D �ӼA���b�����F���a��/]p�)n$]�� ��s���H.oR���)��I�ab%$�XY��FHA}t���UD"��}��#����Ƿ����V��6���,���>M��4����\g5Z~	�����b��.)�^�u��C�e���9�|�c�ھ$	����K~�5�?\DRb�Ux_�_L�\��<k8#ҭz?�����g���q'$��UZ5�֊��f\{��YV�Ҡ���+��zA�kW{w'��8� ������I�.J�1_��x����Rb��6�ŝ���5P���<�c��c�I�lx��YA���8
A	��}孮����� -���K����<����������ڸM4�a�ĝ��GU���2.'�'-���6Z%�5뷘���u���m:?Ɋ9��T��M��}�U�k��)���'��� ����>v�Y?�V/\=[K����k��/sؖ�����áR
H�x1*���W6��uHV&�~�gF�(=%d�V�B��ֱy,QM�z�lܬ�@�3�W^>#��-Ց����,d��*���1�޾�ϲ¦nC<�kG<4���g_���Fٻ��7��`ߢj�=�r'��;��ӓ�54�}:�}*�'���!��j:�O�u~��{V��Z���^��lF#���&Xl6H�t���vJG
�2}��]2�E��k�qo���.�;��+2�1t�ZJM���9���x�r+�k� �߶NJ��G����k/ ���%S�_�p�=L`���
�k�TE!t\ZQ�5���X����Ԧ'�(JE��9`B��f��g��!V`�����x�5r�Y�����>�{�KK�NɄț��o_���&���+���䋾8���߳�
�0���Tj/�������8ƕTj��X`Ã
�ښ�~��m9��|sx]Z^�bdi�F�;
����鎭~G�O8����ӽ���]� ߫��=d*%�̇�篏;��������·	��7s����'����/�X˻O�M;v^�1�Z�}�>�w���BGNU�o���F�1�'���}�.���P�����0�ȰZ�q9���]|�mq2�"�ۊ�=vi�'��z<2�N�R��	Xtη�JC=����.��g�Xl9�u�����~8��g��S����.�o*E�C\��|�!?,jP�/f@c�(	�d#a]d�g��|d���y�&B� �ȷ�B֎����uNo�k����B��[7~*CJ�D��B�H{�'��B�|s���A�9�}�����������ү��+���8XX	��Jh���N�"�'v���+`X(��6�Z�����7&oL���ar?J�8Y{#��T�����q����c.j4#��<-�Tr]v�U�W�v�y��{�Mc�u�k �j䁢2�; �cT�OFK^(Y�g�c�ߛ[���`UNYߥK�P�zH�~~Oh�؋�l*�Z9�-�W�f٦��l[G����n]E{�ש�ZQ�K_�,j�_�^��&��]s�2@����p�] ��~��\vU��Q�FE�2c��hq*
��4(�B/w�໹�9H�|0�P�_6���/��?vsb~�"ٸ��y�AR�0a]9PT�.'3+K1�,����l�JxYy�+�O/ȏ�M���R������%we\��'��9��KS�{��gj���Q�>P?2�^��.V����̧��c��j��q$G���ݳ����Կ���^K����9,����BD�y�qAv���7(�K��� �F{eN�q���R�ph}�]�Q'�t���Bh8`��/;
��cX0��y�>"�.��/N՞e�n�/�q@P�V{��e���7��pA�Z�|ҏL�Z���
ꖽ���3�����+O���S>�Z{�3�%�@�(�r��Z�%��M9�kR�Ț����X���+�{�� �22�^��)���q�FΧ�z,�7sj�ص���`�flġ�ٻ��3{X�:��`��.)����ݴ��H����sq͏���M��6�����U��)��m���臆��ۨ���k�a��8�)�(u�K���k�+��]q�m����M��'��%���� ��N  [��+n�'���W�q�ĸ�4�n@ᮃ&�����Eb��o�A^��ק��!�:W��$��׫� �7�1sq�Uk��*�0��9Y��5���x�5z"a��+?�zls'��q�$����w�����.����JSd��V��'����^Mml�l6�᝔�\�����K�h����	ӆa �ЬjwӒ�4�J򕁼����I��a�µd����Eq�4�-�-�P�e��z0�WM�i1I#�v��5�R�37�Y��c�Z���,E8��h�t_Ք���������T�����?�6�j�j��sa7�! �aP*�˲�fd����IɷU�/���'��8���^�e�S���]-���$�S�m��ˮ�g����c����EdD%Ϋua���e�]EC�l�0�g�	��)��t0���q�bA<ϨRq��A�~�����s��"+F�[��8�A�����ϝo�o�C���؀������oj���GJ ^Թ9��Y�K^E��$���im��W����g�ie�3KD��m�7;J�K�/�V�y�����}@9ρ�b;+�������[k�B��0�m�ͱ�>�^��|�
v��m��m����v�*��vY��yq߳����l*W竊�F8 ��L��=fdZ���D���Rs��D�GX�:�2�7m�lx�B�UZ���y�m�*
[��"p�`Eq��*�\�p�����o&֤�o��Y6~k�W����5Ql�B�� r��*�u�������|o�˝�}���3��V�C�{�Q:��DZ�;DAɼ�+=	Lw��/{7a�$���s�j�]p�$�C+���z$��l��!C�]�Ўcv 0�7<X��e�s��Rx��I��f£��G%~���{/C,u��2���cfw�v�ÛSW�Sր�H��I���{��!��������s9a���[$p����gcs�=6Q��4A��}��JY���~�C�K�^<�/�j�[��o�W�?}�S{/�%���ݭ:�����,����,������|RU��@�)/�B����x������@�(e�Z��2�ɝ�%Rټ�����y�������'W��?�l��ڭ�i.�˼��������g�Ӯ=����aP1���Y:����711�����jU�L�Q��3ts�-=�>�M�N[�H��� W3��`���t L��4��7�ha��w��R誝��Gj�Ugٽ߸� /RZ�������$��B$�w�Ϋ`^-eW��0[�#)�rI5���:�'��PĒ�/,h�2��?��m(С��"�H������2Q�/�?/(+�$�ϤqgmT��ZO��[d 4�����ko��?CI�5k9��k�����>U#�m`��0���)x���֜m�����˲�wcu��o����B���a�f�x*v�:r��l�x8ܶ��k9"$�]��d��>�z[�����d��ɏ:sk�%.�MDn)?L��_]��C�)�%x���e#��$?�Z��=�覸o(Uk��#Vrx���'q��I�sf+0�>�,�PQ���NK�U�s=�Yz�G�I!���m�� �2b�Bu��!^{-h�����RG_E;�ƛ�~��'V��rL��+��"ǅ�B�Z��7�����ve���{-���U�TL�踄<C����=q�5�d�o�wCʀ���	X�
��?M�{;�e��G&U�惌�lt»,K�(���ۜ���O�.ǿ��=�%�e���)Z��6�ȗ�AE��ל��Mҧ�4�eө�ʊK�Z���"G�&7V��Ulp-�VK?>��6�a 1�&=��W�tGi_JN�J�8�*���h����{�[����Z�{��h�gKs.���9�����M�7���t��Ǻ�"A�s��<�>�# �����f���>2�e��}ѐ��]�3s�zf�!45���hk��}�ev��=���%9-2�����7����t=����
�]�s��7�y��A�C��� nR��+y�����T��'���?��^�گ�\����G\��}e��r��:/������'���?^�UG'�W���8��!L�Dȭm�r��7"h��yϽ��"����1G�S�m��ַAJZɽ�5�*�ҏ��x��2?����;��6��?������d��#����̥��N��#o��ULÒ�I���e��=�l �}�7��cxE��Y'U�D-7��ȑ�ܹ���#i��huE���3�o.C�m5$:W&6� ��`�FǄ�7g�;o&�~߻�g����#�nu1g1��9��׳�óf\-Q���ZS�-�O�(��I��r�$ɶ&״#�����G�-�O��h�i~�d�q��u������U�&eC�:(�PU�����
�7��h�=����jfi�A�R6��w����"�Ŏ@����� ������w���hj��~	�`]{V�����fY���P;Ho�(�MD���^�y����x���E��L�ܐ��S[�g⣀U��c�%��I�QOP��.��� �t$X���J�~a�Ns�_��ecv�%9��4?����9�B=�L�Y���NwG ܬ�Ś���6�U���?)SYA�W�W�t��Z��4���,TrHV�67��2Ә���+�w*�b�|I���dt��O핲(��@π���IoH�j�s�"��=vsp���i����D��-�����(�e s���	70�LLҹ�a���q�yc���G�j�j�l���&�X��xڟ�O�mU�w�-���^ �y��"_�(?�ęUH���TT)��SB�NDa�����!�ę����CBX�!�?�K5�Y��)�"�|iQ�E8&e���a�<���꜅3u��'�Æa��Vw�=��4�gY��yY� \����Ŋ6�7��☛�튡�U�r�V����ꍼ���U�[ƀyC��Q2�Ռ��װFK�#�}+- ���ꨠ�V�&(Em�^�\�y�����pSy� .��P���o�y"��ߕD��J��)vP�#� q?��=�Swh���%�xɬ������"���u����O�?�Og�V���ٔWEI�p���c�6���ۥ��Z_`�X��+�����Q�����T�s�ԟ�u�e�#i�����"z
���� *Y+8���!:���EBG��)����y\.��{�-��r�*M/!X���'ͮ=�r��Wl�Y�=D�_؎idv ��9����+�T�g��d_^�<��K�뿰?)f��\�|�ڣ���4{0%Q�$�'P�θ��ۏscVs�~~��n!HZ���q$@��1:T������2ETM��}���l�P�2H�Y~�[d�I$����>�H��1��'Z�G���>��L@�D��\�H�'��U�`g��IVWv�\ �`f�eѴg�\�qy����N������ழ%��W�U�%����5+X/���"v�_�iM��\�8�%�v7{������V����n�����I���y�E��h�^'�epy���@K^/�x|��w�}_�j��4�O��<�����4��T���&�˽)Y���$�����5͹��ʸ>qG(��L�.��5]�z�+z��Y=�Ƚh�ݪ�O���������E(kM�������p�X����Y�1�{bU:��d��D�m<=w�b�$��^=�S1OeN0E��^�����ܝu�K�m)H(���e&Kq� <_p����s�}Rp����߀{�Ҭ�P�{ں�eMn���rH�B�[c[	Yaq�Y��ˮ�n�}Pk����p�����>t`�v'?��[b����b��5�X�ښ+�n?-T�8싏��N�/��ϝ�|E���y~`����/�����i9��L�u���!,�ݶ����{��� �ԅŷ�V/����X+����oc��"��*Zp�$�i�f����Rr��^�Ҙ�U��I�ԯnː��8w9>c5=�댿f���aa�F���E2\��mʞz�yҶ�'`�*'�,�-���ES����=�~:r/,��0��m��zA 5��K	�p��5լ��H����Is.�nV���U�o5����)���l)�[�:����CR:�$u��y�j�ww���ٍ߆YiL/h,X��P���إs%=�H/�%"�0��W�v+_��|j���q��?�NQb�q���a��O��q^S��Gs-_Z,��*v5��mWD��N���FrAoM���|5�<�s�U�-�\����V��3]�V_�Ψ��}M܅�Cp�k���pcT,6ϨB�|�� �gO����ڦ�����J���C�$�������Q=wn�`1�ӆ誁z˰�}]����
	O������h0Q����	}/�M��*0[�����ǭ���(;��~ů��P	#�h�2)U��~���%�$�:̕�[e�G�S��U�z[.�IH��,�`�vdl1�.�yw�#E[�Bt� ��;�~�������6Yݸ�ŷN>���6�Ycð�s9_Ώߟt�^/Ո`��'�2_c�~�~�����=����)��<L�_����G����
Aq)љ4���^�!�!|N��qSx�"hl�)0˙~+Qb�f�!��١��NʑXW�6G�@LW��%��V�l ��}!C���Wi.��
��MtĊAl�a�ڱE��?/	�x� �LP���?�@�{߅�[��z��z<�8��N����ߒ,��)����T-����.�������}��h�luo�C1����K�ɼ䠩@'����D�m8S��z��Q�M���'�_�����K�Ћ4�J�Xq�h�qc���Տa>g�]U�'����V��C@���K�We�jأ��g��/���[iN���8�+1����*����[���Lb/��%"��o�V~�%|��Kv�Z�+�j����Վ:p�;26��#�*�t�U�h�)a��:E:��^\����O��[�;F��뢽��R}*d���/�XY\��琦z�&��D܋#ɘ���FL��J�>�N*�r3;,�����p�&����v��{���
m�m���Z�O&|Co>¯�M��$JY}��b���4�^ڑ��;XNc�����#�Qf͟}����:��]�0���ӣ�'��K���%JT�@d� ÔwO���� %�+&�T;��Ì�
�7�͸�F�ئs��/��o������C�L�a��rÛf!z .�V	��p���ʒ�T۝q0���d� ^9
P!g]B:�H!��9�w٩D0���ɔ�F�S���~gx[�w��$���RIP�/� x羁m���� �B�W�(�k�(]!U="Y�� �s�|g�*hwynܯ�|�vqy"r�M�K�E��A��Xvʔ�o���'R��b�@��+|1�s���X���wNQ�jM�G�$j��σ�Zv����^ϻ�2Ӏ��r�0��_�_�~��آ�-��N�kY/;�^Ԯ�R:��'���6h����(2Z�"��	�2핊�qi�_�=���>U�������tŪMx�T=.��)!�5$~��Eز�J)�Ŀ�"�I�ؽ�!�>�D��팗���y�Q<#ܺ�a
s�y�;�G��{0�"Cd޻\<nz}A��gw��\V��@��k�7��Vw��T?�+l2&���&�����b�.��gL�!=���f�)l9�i��`�Wj\g�^����!��.vlY�E�rI�}����+�Z���;�

�j˨�G�{e=hƄCO�N���PmV#%�̈́~���z��L$�{D�h?Fo��C��o]t:�J���nT��/�S�?��/���IX&�g=Y�q��������WD�g%�!��SE�I�4n��]��{������$�-aX�j���Raj��-�,��7�=�M����/!�����߳���RCb��.훑Gp����ڼj�pZ"=<�����,$���X%`Sx>��,��J%��tI�Jk�jOA�*�+�a��~��������I�g2.V�������"��Y(|��G��YX�1�Y$��6%�� �ᘘP)���wD��,I���s)���t�	zy���X}�k�t2�����v�#����}
����c�\�7к�$�؋�������P�]�.�k��_���n�/���Ɔ4��n4��@�}c��Ξ|�B��Ȑ�\�6�W7�C�� Yݏ�YV�P*��.(5�=([����� �*�Z��R}��F��M�
�fR�o�YrU�T�d��*.��č�Y�ώU�Ba����7MM0M9{�&������߅�_0Ξ���z���ͬP~A�S�@n���Ѝi(��0�#��͚�38W����������^��x��M�}96<C�&���̿��u�R��s��v�bl�=��Ci8����<Y�����_������Ҳ֪�H������9�PI��_]��	U�P3������#�bd��;ل�0�U�vZ+�y�`\��"s�+�:��\� ?M�/;��g�}��uj�?�J�����	c�o[�6�����Rݓذc��g��#'��ZVCD�5�������z��w�\xT7��G��֮���g�
��D4i���^f�y�_��1�m��+S}��O��ď�u��ͣA}�>��"�&����_���$��M���6��q߳#��>����o��ڿ��b�%��S�Ѥ���L���ي�#د�R}r���H��x�k�턝'�2c���X��zY�o|��G�o��H}qʱ7�)���_
�<�hdl}��kr�݁m��U��9u�g�r}˜�aՏ�
k�Y��$�;��~�UtK�Vo�~�n��Brx�E���Vw=r�<�#�=^I�c��|�](C���d��!��k��"���FnKw��CDUh�J٭�q[���'c-�~%���}�5��1�P�WZ�Mg}��d~�O��z>���#{{;+�Dɠ��q��w�������C��R�Yd��v����>E�c�c������H�}�Ǉ�|KZ�yv���>}.E'K��.c�T�J�[��>u�)@E�<�����O�\�-���o?M��g"�}��p��et��R���nX�!�Đ��;�Sh>�+]�x�ق��)��%w�iS����k.��g�-Sf�T�`#��l��,�vH�o�o�"��%�2��eI�ؐW�N��P�0�F��gC�щ^���̋�*�,>�Q�Y�$�
x�[ϐS��x��6��|�:�'�L���j?�L��.�i�j=y͠$=}�

b|��Wo®kVu�q}��P���~h\�2�-��B��4Mt�65TR�&�9yg^�,��J��������s2�WR�k~�|�ƾ�bxl#�ϋ�w�>fe�r��e} $���3O��uR�P���W8o��r��^��~-U�)�t�Ѻ�7Co���� �F��Y�0�v��oQ\�À��J���\'`���F�l����_�BgY���%s*g^֪lWgW�ífW��$�ʖNasZ���N���a��Q��.��y%�[�Mf~C�9�LG4���z!k��o$�2ha�>�D�����H��]�������^,_&S��ƣu?z���ڭ�_������l>y���ɬ����y����_qm�c���ɝ	��Ӽ+���|��z3&�N(QʴIL_�?E#�BD�O�AX@T2~�*l�\���P��׮&��5��DKQ�#� ��ӓ�7|P5���dc��؋�a�P��'O\E�yą��9[f1�8��)E�9�s�Ǡ���>�4��M��m�l�rì�C�&���n=ٲ}^���S���D���Z�O�u�82��_����
?�������C�^��|�2O�U��Aj���ѣ������M~��Ƕc��w�j���	x������6�:�X�3�^B�4�I	�4�F��K{�a��9���_1�$�(�%�t�a�|g��-��/���4Q\C^�]����h̫<�����R)騬gG:�������v��-?C_�b��U]��t2�3km��Q�.�%��)�Se.}׊�Ͳ�%Z}��ǲ�䮡,wZ|g�14����Xe���Ϗ�}�ܵ��v��+�|��w�d���9�+	�x��p\���t��2:xl�ְ�����7��UZ��V
�����Z?Ʌg$�(�$�Մ
�ց�hb�鄪�ԇ�M6��Ұ����%�݂��Í+�4��������Oߡ�U�����g8x��X��M8M����'ѯ{��b/,�7����'��y}�2+�\��@h`$��m%�d���Z��_|�v�5D�9{������\@��e�ݦ~gq� B��D<t�c����%�^{r���zRCC*��|�N�{�ɜ�J�p,����y.�y���'u��B]V?C��uc[� 397���&,:�����{~���c$w����!��^:|��~i�J���R�UC��]Yʇ[WdMȇ%�MڮG)�O��v>���|(*EMzv��*��
����O��f�Z����P�xo�3�WE��mC�Ry>;ޚ}*���a�y�ʧ~�@U5r�|�	d�k�P���g���v+1�o��OP�MC�a��3)�5.�;���J+�g�`�����.�/�!O�q��f)%9,m�{Y��/����=%r��<��-p}Z��}�Ta��E�^K�m�A�����e�޲T��]��y�VZ��e1gf���� ���h�I���`�|ڐ/�ҽs���v��h�"_t���&��� �"��cE��`���u�����NM֦ͧQ��ĉ�/�y�į�����3��B�zA6��#��#W�ޅ<Ȣ�/53��;�e L����78V�}7J����E��iO��t]˞A��Uxr�.�M�e0�k�[��ŝ��o�O�H~�F��ߋ�E�?���f}U�\D���f]I騌�f�$�ټ�r/Q)?�9mB�)�J��#�7����x��]���vbX��{8����^���'Pܻ2�{�j�7y�E�@���.VUC��tm�6?�������t��j��䇍.���2B�c�Z^��Sxø���R2�����$[>�#��r��W6���q�3����Ӳ)e���i 9���_� Cִ���.�H+B�)�c�K�~" .]��|��#�c�fiv�!����+)����Jd1߃d	�,%\��r������#��������m$��Ip�qH牬���H�q�E�i�<������K�K�:�虸��g����a^�Ņ��%�b/�?:NU�h�ݧw������U�Y��j��N$��e�w�/���ֱ���Vt"��O;3.W)�R��>c1aq<�3�^=�vE�AN׬ѕ
�^`�/���2Bf�	v�9$���-R������WHQ��J^O�e�s,8��9g{�$�.W�|��zXNV	���
N�+�:!l1���@Q�VC6L브�t��Ġ-�&6;����z:�_	���͍�-ux|1v��~��:���%��\�1P�@@nx�L����Qi�ak�|e!�X'�O������!�&�\˻\��kr�(J�E�Z��E��=ԃ_�_^H�Z=m�7����[����0�@��15`V)����m$��Ij�I�l��0�S��+��gE��]
d� \|�0�8
��� �zc	
m��<�͉��a�<zх����X�=�{����z<�������}%���ş�3��^�E��Y��|$��w���tL�s�]�)�	�~ps�9r��)��f��׮��aE��K��̩�fra[��2��Ϩ�[߷��a�b$�=ŲV�����3{i�7}�=�����ڟb�C ��#����1f���E<�>�>S�\�JQc.�t�Ӧ�ŪO��V�S�bl��;�o;&��.�\:^:E�Hcc��)hnPָ�T�>�r��=-r(��e�� Q�cB���H�k�p�P�i�UcL9��K�w#zS�K�_� ��T�eg,,՛z'�ej4� Txe ������Dw"<�7��3�%'_� `n�����hy�Hg�xe���i����c�aΊ�8VO�e�m����ȁ�#��?6��Ke{�h}J��. Wy�������bL���8顖����t.ꕟ&�e��
� ᥚ�a��i�����)�
�(�j�cO�۳���N.S<�m�32n�l�)�0�o�JͶZmtx��Z���t�ֿ����,)���t\�����C��'%��(�&�2�������ң�67����]W�ޓ�mtJ)�st24I:�7p�7kLdk��t$������R�"�l��x~{,�����?���d���/>�M>v��x?��%���?��C߶\/�B7O���+�f������oX��w�R9�y����:�Oרq��l4˻f@�b����qE�~���zy����F���������<�G����J����J��������ր4��C�k2T��/̽+~��a�Z��ͥ��<��0�� r�P���R�zl���U��.w��&��U#(">q��+�[�Mś�b|=(��h�)�%Ҫ3���	!�L��[�UMQbq������	��7~�:�^���~��o/ B����<��7�%��f!��5��������� ���1�wv��O|}�$� �Wץ�b�7�!���Uy��{�'�R1�&����)����EC�8c�����ݻ��j��e���wDRT)�8�X7":sQ}Ku�m�bk)���h
~O�I!�C�Y���7���ϴ|������T�:��.s�Г��*o�������{�~��9c5�}�bS����~s��ϘT��]| j$ށ�u����K��Jw���gÛŦ[O�H�v�Y4ލ�M��ƞ�������XԴ�%�L��xs��7��h��~�������2]E�sб���H�����<�ZP��z��ڃ#�;XQ��Mm>�0�nʾ|"�UO$(��j�>�1�n�~<{3������[���o����E��/�(�j�����}��̤1���	#2���0D}�PuzW���dӶ���͔m�`�L��l�`]�`]kgBi�ħ΄O��/�܊�\�n)�(����I�~�ǈƨA����ќ>����ur�ێ�ے9j�^���a�����q��R@Ӛ���gؗIx-�:]ERr�D�"��o�����5~L��*�]\����;�j���rfMe�:/9�����$�y=8���A��L���@SW��}r�(�;�Vо)�LC_���bhZݨ<i*a-!@9A4yỆ���n��E��6E��Eܟ��\8P� �bB;��\��+J�u�������ϯ)��~o�./���n�����q�`��e!R�7q0J���J�>���b��)���1p�˙
k�.�$j�;ܚv6�#�#δ��8��A�V�~_V�j��9KЏ�fo.�����]-���Y=�����·�@���@t]X�)Nd�UO��+���k��"U��|'=�"o[�쌭��� z��8s�yZ,�,�2K�Z.��!bU�v��G�J��\��~3^��6�v���� ݦCe�8��d��|��,�ܱ1�}��V�16:uJ ɋ���R3\ڼ��� �T�k*��#�r/��un�f>�������q�z���K����떦*[X��.+�Td3g�QM��-�ι����F�A)���*b�s܀^[�Yr�[�� R���4JG��jȧ����V3�rBśf���iF">"xWN(3��FJL��� S�F>��p��Rv�X�--��}���z	�E�1�������M�!�J���A�d�r
Hf�&ᜱFn�<�Ov��+�eNCs��u.���F��7U��d	`��	�ciE���3�ܵ��θ�_2�(~ù7�V�ث�T��یÂf�����y�L�o�q�~s������2b�C��S߼�2��Qm���r�I��B"��*����j�6�>�`���3��+�#�������y�Ͼ]r�S,�mln�7�qҞ�QO+D">�s^���1���7=��&���Rۼ,exE�0���`+s��]��0�L�B�~k+)ٳ?C�,.(����y�G)J�	m�z�������ە�c_��a�ةF{�:;�ՠ�ɯ�Z�B��˅%����T��
O�' R�{^�O�	�}�|��c�kn�jP��=���=]��3Zo�є�ٛ����-ʭղ,���Q�n����h,\^-;�b���{R/N��e�t� 6(I���jr{x��4S7�hRS��R���ЍĒ��P��n�f��`�d�I�W^,E�Yoz�'Ku�W��Jy0V��̇���Z0W�ɸ�6�Z��h�&`�2?���\��fɾ�iO؆H�J��K�ZrT��Έ����g�$3��ʅq���A�������?���j0wSxQ]�e��j.a���$�8�QSVZ1�쌟�6O�o�����η�)�)Ta%�&!&Q�~�w(���]E�[���FVR�����i��g�!�O;�.Ց�+�C1q�L��yV>�@���&�Q�>^��A���DS��-+��Ɨ��փ׊}֞m_�4�����l[��8ܧ6$,�A��R�K����$��,n��/f_x3m�-�2�هx�c$|&*��_q�	7'7�Υժ�Q*Ӏş��@����(�?7_�O�����>��K��}H(u��&H+y��T|���z���� �sOſ��o����5�Ui^48o��r޲���l1�<+vt�/���V�؉������/G6m.���\$�튌�b��H�;�2�_�.��@u�X�_������,]���.m�Ӫ���Q��,���Y���tH����u�'[��-�'U잏QC#W{wD�kO��6�L�j���4��e~oK�|��0q��=� ��(����Ϭ��$Is�M����_�h�/���#`zG�� wgs��������Bt�]>�"�������Tf3�h:�
�� 1�fx�o~��%4�7g@���Ԑ4y�L :Ϲ�T�WW��q���Q�c�T��ь��D�)��G��b�����|Rc)1J�ч�^��Xm�	�&�6'��@;��*��i�����P%miŐ��7p�A�4�)������=p�b�e(A��	իJ� ��� F���Oq7wk3���} �Xm�T��j�=�s�#&b㧼��7����.W�c$H"�r1��;#�s�c���̷G[������ס�۱V�j�U�/3b�jԣB�.�o~��K !� B~���ʤ_Z]�k;*���-f��#�wV���ۇ��A�vw�~t;:T�LX/�U�a� ���������qj��Y�Re��H\k�+%��^.�6\�θdj�e{,���)�a��n(N�7�#A�W|&�S����̞�˫!���&c ��|jwqCP��%�E2Ѯ.Zn{&fV<6���,���I1�f�S��|�dcёfR����^�U��.C3�v�Q	�r(����++�:v��Z��NҀ��È_�H�ʚ��`h�(}�U��O�	���i6O��T�B�$��l�+�8�L�?�=.Nv�i�����@�,����{�J���W0�I�C~7I-�J�m����{�H�f�1�Q+���o�[h�}��a�;~X��'��I�X��7��x�OR/���P���p�#�+�&xz�_FϢ�gC�/$U���V&;�q>Y�m��G~1��z=�PHb􊪖ߣx�f�\\�6���}����h�k:W��WRu&{ E��,�L�P�BJG��Z-w)و�����	yH^~7o9T`���0�FRǑ�&������^�Ayw��Ҹ��n�3�����uhJb�7��lNKw���[�z	�J}�r��e�����w'��;/`[YXMnt]�\���;��X��=1f����{ؿ˚�6�5u9�	��)_!���L3�uF�ܟb�E�B���9��.�Ec����E*��=��.�cx�7hk�9�z%��a�]��<�ŭ�w���=�Nw�؎���6q+بx�՛z'JR=�D� 7T�X�.4����E�KcҒv�<����| ��	o��צ�:�2j�f�4�]k�N~���F��$��Xr�i�`�a�c˲��D=N]�ߎߗoT��i�ȴ9�4]uT�[�G���Wa@�[j(�n�i�zD����n�.)i�n�b�����~����>{��s�8�L�?��ն��Ou��ԣ�Ӳ!�
����ĕ�3��9ᵹx4S
w��d˸ִ��6�Typ
ù{��֛xu�U����D%/2�<=K��a/�P���XsM�,���,��.��#,�G�.kkm�����\�.=o����Ħ�+�/�?�k/��
��<s�p�ͩ��Q�:)� ��
�g�E~�"���q>1y\4X�l�4�]���&6�}b���kY�9�i��| �T��@^%��d�:�ɢO���őSk�%}T��vm�� ]�`�ĒcC��qW{�# �޶�Hh\
X%5ݛ.�f�L��?�qJ���A�j��.g��& ^��^�m*:�܎��iz0yv��!�)���� ������{0�,
���l��{ ���*���$���4�j������2�=��ǴL�I�%�Mn��m-5/�߮[62љ��O��O�.����[0ػY3l��N(@$�5)�R���fJ�N�����v �㺜�o�r�X�UU�/Jv�p�\W!�o����I�M�RiF�'	r*	%�ƹ�Mq�u��Sl���sz���<FK���Z2w�STR�]��J�Te-��
��u�6�՚��Si�Mn�mn�5�2�9�	���@�u�Y��u�2����Q_���XL�N��?Z�w�1#ں��|�"jUb@��^u��݉��֓*�>1����Hc}n���V,1(�)�b��A��\�Y�Q�4���+�c�VD����߸!)��Т�|o>e�}�Ձ�0'>�<�V��+j�QS���8.����:�5{-�qġx$�]\#�H�NBt��W�O�f^xpW��e����`u��:�_OjDEG�G�0_ԇ�#�1
�h-+���2�Z=&bXl��kp� 2~5�8�|��A�L��;`�	i���:{W7��0,:�QMcy�!�w�Ux� Q v��g�WdP��]�\�o)[��f;��_�F~�0��L)�k4�>�����v�?"y�����s`�g�FVՅ�-W�!lSs%3��6t�#;��òF֫1X?�׊M�f]9\V�Y�c��M>����>��Ͻ&�sG����j:��2�LZȾh�Q\U2̢$I@�[|Y4S<7���^��<����0�"1۴��P�e�{��E���*�*�X�����ֵdG�	~T?�ʦ�es[���,���QC�G9|��T��OF���z��*(���@�z��y�1�K��JV�f����}M���aq�u�����s����K~�S��u��tQ��N�#p�`�ꊍ������֬�ƬH�Q���ܫV�5q];����2�}r�)5-Gp�Ǟ2�Fث����WiW[��v\[{n����!cW��ne-kQ&�^�l�&ҭu�s��ð�E����U\�n{��,3�t��"�L.�Ȧcd����u׊�<{���<!��i�l{�E�;δԷ�B��?����EPR��i%���X;���~S��m�.�����B�6��E���L�V P��H,�x �#��A]t��Ia�amK����Q=�R�`��U6�S��N����N2�0ٺn��~�������\�]|��ď�Kl�Մp�A"5$��.Iof��'�R\�F��+w�6��ɓGbڵl�����P����it�n"��Y���dvq�p�9^+1g�4������{��X���:�Z����M
�ޑ�P�?�ݸ�j��Iv'$�ݮB����&�%�k��|��GLVt8M�=&V���Dz��68#
Xu`1~��}��b��`!���=�k�'QF�gF�[LU�/��NH�f2��c�?n���n��|]��Zp�_Xc�I{� {�Xf�K�9�x�_)��;4y�M.lk�e��RT�J,�����Xq��`͛;�O�&�U��*��d�}�?:�PY��/Fw�q��,0sK�a��6Y��N�WT;׌��i�:������磑i�GSgA�w��u�zfX���Z	yF	T���qn�f��n��[ �`��{��#f��e~g�mns�)=Q¿ ����UJ��iy����b �#�S�{�5B��ב/�K�b<�#��N3'PpY��|��^�����էX�?������R�1!\�e�?8��[�ãUD�7�C#�9��N�<r>��g�8����	��m�M�;�^��;4�KW�����t^G�����B�9��-[ܑ���BX�7
���u@H��\��u76�3\^���zh���o9+ٹ�ڸjՅ�w	7�{@8̾��~�g�U|r�kW�t+��6��i�k||ԥ��yQl�*3'�i+H�8x��w+m%�����:����!�7�K�v}�o���3N ���[=��L��Xr��*q���D�B�w9Lkx1&��rZ�����-�Y�G}+�)��!��X�5��Ĕn
��-����M������|=؊B�Q@�ݣ�t'�g��c�n��*��G�@�L2q�2x���UZ�H����>I�#>nmS��@����X�y�K���Ψ����I�wף,ԍ`�@50�M�3�i���I�l��-�K�@�4O�_[�>���	ި� M3����~��`�e���X�f�P�i���y��R�7ЌJ*�nb JM��D��:	<�~=@�R|�je�X0����� ze����-Z@�2��H1��2}�H*�������O�f��b���Vi;�h�-ǧ����G��h�dD�����5�����e�)hYG���)�p���cU�@����=�M��RQ���h�O�z����դ��ë��R;��_sl��:fZ"�DB�7������@�`SK����M�_���
;���'��]TG����2LQ����3�G���Op�65a	��'O��ܹ��O���L����M^�<9��q�τ���V߽V��kɕ�����aF�V�������*4IR$�İ!�;�m� }��f�;�Ԡ�R�LEbB����1._K>LB�>�b�]�>��T���N|x��w9��b�MR�Y�t�_'��ׯ��߻�{�{���_5���k�VWM����4r�J��jqS3�ȫ��mhK��&涤9J�qh��e���e�	�FFםS�����)�C9�\���=G���R����O��S��5��[�i����U��'Xx�z"�#���'�.kl������q>���Ա�tN��^��0�^�Xu9�9	<r�2}�Q/��^.F�0�^���aBq�̒>��~�+Y�/C50�X���^w�Y���ZF٥���<�ux��es�����^�~��Rn�ԍ�����%��O`!���	�C�`u���mĊ�;����� z|�����h؞�Q��m7������d�>if�.D?q��P��_Vg%�ї����L���w�W����T}9 ���rem؟>�s9)[[4���T��!F5��f$�D�!�Lq�E����kb��(�lM�@q[�Y�:y�X��!��Q�HӠq�7P����1�������߾�����:;g~=���=	&�������1�޶m���:=B�a�*���0q���.��/c|d!,�?�$���u�t��;˖�bE�vh
���OP�Nk����~^������D�Ҟ뀼�:QM�yn�l�����������n�t�C���G7�T��0�7�&d�4/;'��Q{duqj(�{�2=�`+��E-��
{äM_��g��t��u��MYsMn^���q�8��C�w��9��#��xU�j�nJ+�G�S�	>��D(��֗`˼��]��5:T���>S=�#����z+�k�-8�=]�Ⱦ(�[�I@���7�Wa�$�u��R��+�y�r��^�A�'�dPeٖ>r����Y]ZF�)�{ݬc4�v��5ݱծ�D���1Z��v�L���8����2�^���Y��#�(>w�L��u��_К�<3�0�d����c��������-��J mv���	��u�j��r��vb�-�;[�:A��&���n`��'hD��o�:m�w԰Â�v�tȫ�lKt�{���+�S	4��p<����9�{5��?0��<��Ct�K���M'uΣ�rI����r5(J��!���3�����F@��,�?�'L���Q�#A]��I�,��6X���^)�W�����%���ߌU�����	*�E!ĉ���K�6o�!�3r�	oM�ܯ�aE�_�C� CA�X������	�Z�:���}������v�7�xWy}��$A]��=�>�<���7I�4��b}`ޭ����ȱ�oßfn��u���ү&�TE��[�ɿT��[ǅ�\.��ه��whᨭ:]��Ձ���^���h�b��0��o�����]�3;@��˜�uU��c�������l�]�'5m��DЦRǋ`�~�r�k��ճ���v �|��f�Z����z�W��>=�����>��
N�gS ��n��M/��#;��"NE��y����/����\\c��sZ�?<��f�?����KȠ>�C��R"kr2��^ܓ���f��[=��7�A"}�<�N�iޡ1����.�[����Ab�_Ի��7!��`�fj��Ѳd'���Wp0?��Q������Y��ٵ!cwi�#kMM����-�K�{�d�����Y�1%V5L�ȉMsޤ��� ��i�-(�W�Ӎ�=�GND(}mvV�I���^�߅�\�N�t�%��T�G*J�G��oe,�s"�+0r��y>�d�U��� 5��J��Ò%է�.~��6��ƙ�WߕMr��W�o�9��R����O��g��e����s�������>�I�Fq�?6��U�|.۝3͘oB��l��dk^����sR!k��vK��4A��
_{���'-+��J��r�k�qS�`��9��f�u{#\�VV���@v��0��{׸���4�O;ФQN�  �&���@�V݀5U-��r�4����\S��?�6\U@HaCwb֖�Q�sr�X��:�|0V�N�*l%حi#��-���z�߮g@к�S�D���/N泶�ٲdU�z�:Au(���(R�9�6����k�tcZ3�����m��Uy����'��U�+�?�	�	��I��3�Z5��
�t`p�r�$
e��;���7^W���Y�z�v�8������D�-!���۶��,�3���m̚��A����Hw���[����7�6�u��}:ͫ1��U�"U�Ȑ�"O��Ӟgx>����H(��jx���y����ٽ4\tªh/�D���M��������OWfV\fz�.��.�Sir�Q�o�x�c:&4��僿^��JUuC�|WC�����f�bx�c!s{�X��m���Ġx��m侘Ԉ���9r����p���<ƿ���b���(�
��Yi����S�����M����s�(�h;��s�i&6!�g��J�	mŚ�_�S�Jq���  �[Ti���`	�zHb�����/]gl�����}����o\��6���O����-�=$}�~�&X��&h;�J�x�a6L���+�l�-�7f�C�}8X������E����9V�E[�o�͵-ZI!G
� C�ri��)�%=��g�NY�c_����(�_&���ąuK\[Zё�G7z(���l1/�MD��6���O	��QL���<��/��Q����P���?�r^���%"�,���k�n��e����T�,Ǯ��Y#�-�/��O>��X�������f"��Ѽ�ˡe�c�N�b�5���詖!�	�����ΰ�j�2}��n�Y��^da����}>Zՙ��n�B��-?.�M�~p�j8���0���'��\��>� Lc	H�ߥM�k=pC���eb�?72`�ݡs՞��3��:���|'d���610���e��e��$1�dO7��]p�4,�X`�?u�SB�1�̗y��I2<u�� �$L{c�r,����ݧ�����?����g	���}�(U�O|��o܍0bzǗ�X��1 ��5c���+�C��"��y`��Ud�y�Q���uK9��i��E
4cV��-����u�%�����n�E����δ�ؖ�̀����5 �ц��K
k�,Hm�v�,90.�� )���k^��1�{'z
o���m�Ĉ�U��ڝ�E,�
f� ��Ai\���v�J/M�y�fR����<n�;�>-��	W�`. ޯV�r����c��-�b'��]����c���N�%��E���U�ٷ3t6[�\�����@^�������f˘o3�M�bz��m����S�yrX����/1(-Sl+��c�/K�!H��X�����T1%�I(�NB���-/�ǐ�^6I��^�����v.Jli���Fn�xpS�zQ+Y�Q����M
�-Ŕ�+=��eIF�(�<��@��@�+{�F�;�����&!�vKh�B*5�������*#8|8e���i�:�*��z5�����v�������,�|�Z���6<���j�>'�m]+cڊЊ�� Ȁ��c5@����)�^�������f�ʟFO���U�� ��J�
i�
�\��
>B��k��-~a2Y�V���4�V�lQ_j������h.1��g����K� �qbF����l�h�����F��~��̋�vOi�x�y��2=�X�S�e�;u\�,�vb8!|�۳ X����e=u�y��l�d����f���Qn��#�u��iI��o����zo�5������.䪒+��
(ݤ�����W�8�3X7 ���?W�LJy��bh�K�K�yl#_�/? ��s�x��m�f�ήIʝ�zuW:Ќ@/L�����w���7���{���|i��B��� IS!Tkp��@j��G*��B�Q���!�h�@Y�n�sp	����~�����<����7U�Q�X��&�<t��p�|_�|�$���������7Y?���\���tq*�Ck�'�6,w[Oxz~6���-�S���m��?��M⽲�z���N��v��,9�8�Y�#�pc� ���j�MaB��˺�Ea~��RѤ�6�1ۺ��+�!�R,}9�W��Q6�b����:3S�gׅ�Q�Ħun>d�᳿b�-���m��(���a��&[�h��{u�|�iu�r&NI�m2����M%%*�^�Y��U��$�RXZ��L��믦�Lۚ�X�Hs w!	����$�y��n#I��������?�yn�U�UY淎ZM�n�0GݯE����(*�1q)|��E9��_%)=�Nh���c�0��t7��������0[Ѹ��+��:0���/�`����ca��Cg���9����q9��5��Z�i>���6r��2H:@! a�~��#)Ҿ�}��-��7
��չ7��x�ֆB�½������TN �{TK+�����t�Y�S�2��c����7��9cƭU�B\��v��LW�h|�]ow���y
�b.������i�$s���!�e����k�ߒyew�@���s���' �iCa��$͖�_J���w��f-IW������&Bk3��f�g�KO��Z���Qu}zZ��sI���r?�9W�n��H�Y�A�#�\o�؅f��s;2�*���o��;��7��N@�D@gr`S���+~ Zh\\��סZ�p��Ju^�z��ˊ���i/�I��Ռ��F��@����2V��<
 ���d#z'3����>q@�i�'�����*�ŧ�[�AM���Dl7(�W _/*����&ο����S�V�\1����	�NMպ,�V�����t�`I�3|׎c����Oh���H���� 2V���,�zA��-x$7�1A�AC�:H�*��ǲ�Go�f�&X�T��Y3�E{����U0�>��.�l��M�9��*0��;%דL]���;Ui{b�,���Y�������:m�l
}l^ef�\6�9��*�o+�x;X�V^]/������9�h�}@����R�ю��i�|c�D�
g�+Ͷju[�Ρ�E$>�O^Ͱ�f��a�).�[���ť�+��Q�6�$*\��� ����e�	��y'� fm)08���A�6b�E��	&Q�������88A���(��C��O�v��[���j�zzi����E�jS-�dB+��xx]j�9�F; -H�S?���8�R�}�@���dL�QWl#�vv�#��^Npcz�j��ћ�8//p�,k�+5/ڒpYj~:!��ѹ��)n�i����YW��F�`sݻ��,O?�?Xt����+ϕ�m��_ЮIvJi�eZ�׹��I2�
0�Hv�eCѥ5x��!O�]cK�#�-qٰ�UCI�i%�JAtN-�V������T����v�X��F*[\��uI�Cc:�C�\��G�B��0��&��A����I�yH$�r�>�b�;����aK��,g����IH�4����<��-=��g[�K&qX�wK~�|$3о�E�<^Iiq{w$W��7$N<�Lι�0{��T��i�P��=�	eu:�.i�=�B;?��GL��F�fn�:�e�qM9��X�8'�_�1�j�� o��SFL�3������������s�q�2�agl���"��H���1}�->���>�A��6�
f�i�8��[Zi�F��0	���1��
���o�7i��-�㌼�|��#cyj=S4�½�Aqb��Ŭ�{���_'��|��mYa�m�WW͑���b�'>����yH�j�[��u�`���Ԗ�9�/�>lQW3mY�8����8���`���\��4�6'X�WX9G>ԡp�x���%6f׵	Ȩ���[qѡ��=!Ց�G�x��� ��>�:��˺�SU���Y�5[{�������T��uW�[��,���5���6�MD0�yn3j�z���ʋo��)X�g3k폪]U�(>6�#'A�|1Us���l�|� �%B�F?dT�$�CҾ��(���d܄Di㌏���Fx�q�Ë�J�81鶴����f�%4i-֪5>w&��`O��x3�B��ʧK\kjS�� ��429��Ċ��~���T˃:eT1���H��n��ꃩjO\9�l��b��㤏�iqR[c�=�wd�t�=��S:������mf{�1�(�;�@(ֆqp��&�5�V���ơG�]=E����[�릭�J�e��5Z?G���.|�e�����9Hѝ�9�I脖�؁���(��QQ[�U��w����]̽��=�ȡ�^W
G�(�����đJ�sb�Cw�S��m:�������7�1���b��{�܍ʀ��~-G�#��UJk�b�Ǡ�U7��Zdn:���[�`���swo��Y�R��pp�9l��� ��In����+�Q`m�$w�$��*	�a�E��u�M� Ƣ�������q�X��퍅�>���=��)g�_^�PvR��0z�<b��j�9TH��N���TV��p
��_��h�MB��!u�om���>T�M� ����uL�H�s>�sa��c!�ޚhP��k(`O�����^���Ԏ��t����HX��x"K�����^"ry�ǣ�S��+u���q��O�:�N�wG1+f	6�%8ɹ���L��_��M��W��{�c�(OD}Z��m�����������E,���A�J���㾃|���qJ�KBE�װ^�4���
a�+?����.��?���x2w�	O��vi��h�Ug�tWg��&T�H�d��4���h�}�لO�ϗE~8/(@�U��F��	*��.N{Yjw�k|���]�R��ܽ+��G����J��]�p}�������46�IY<w�\/o����_�O~v�^�RLz���8��nᯡ!˚[Y���3���Wo������y�X�I0�gd"���9�kI�K��p�l�)�����᜼~b���o���A\	nS
�4�i�-��ed�?J!+�d~+6 ��GbO���ͩ����nS���?5���	Zu^��T�D9j\��Ȅ��F��m�&��88'���� �j�+�
Dy"Yq�d�"�7�*���	XS��^2P�}Cr���	�<��P��fh�흵�X��O]�e���8�VsR�Ӵd�?�ջ�	����t$n�&\��G|�;�XY��g�V#i��##yz{/J�����&�<\�~dV�9E��Ǧ�=�vDgO�#l�j��C"f��>fV��0js�m�Z����`V�)�4NF�5C�my�Wqb:����8���Y����rEp4R9�}{j<��:f)�i��j	&�Z9�M��
�ٽ�}�h�&NT|gԂ8Ha�5�����t D�G׮�������e��x^UKK�u,צ�&7�a��=�P��`���b�o�	�yJ��ki��d|�X��K��?-U�Vtzx�JzEuW�Y�1��-�ԋ��_e���,�	�ך~��^߫z�#;�O ��Ϊ����<N��$!9���0�q��x�Y��<
,Y���u�i1���Y��m'����[L��w�u؝�Oɚ*�/I}qwlby6��~t��t�[���c���d�{�i��t��\ԯ�*0�ۢb�[O�/�;�4`[n�ן8gh�ǸU&�JF6��	���tL�Ҵ.�`!�U���tp&��DжJ����7k,��eAX��|'xNz�-�~�m:����^���Wz��d�C�ʛG5�8%�|{p��>���{�N.��a���M�z��A �y��(�]�7�$K��E��K�k����Qu��9|�E#QX3��ձ����U��k�`0��I\.o�O��\G�j��e�(� 5�����dEε)�޹�z_|:Spw�%I�b#��k���UTq�o9K^6Q�+��_�K�󻟸���BWQM�pR@%���\W+����ט��y���+-Z���y�Da�6���uBj�Th�Whes ��[�]��2���8������>ϼa����KTB�\�ќ�D��W��'E�G�z��G���E}�k���r�����_^%z��xy���./<��n��s���.zQ������%~Ȗ�RE7�Ͳ�a��V�
�*�Cy�0����OPNucIm���I/X�:C��3�4SQ�ot��1�!	�>Z�W-��	|�J��C�a�ɮe^X;1+���'RLoCg�=xz)t�"���6��H�l��+ӓ�KK;�^J829�������&�|�'Ͳ�	-�S����><���J���@t�T>�$n�x�^�VKhZ�&p܈��3�j�%��#*y�~�4���K{��'H�=�t� �h�B�;M����4�9�f����u߃�8�.�T��� D8+���ҩ��;5;f=	��.�%VW�%(�b<xɡ�\�������_�i��jp����Vi�*,�D�3ލ�@�uAR�SU{|k�V��Ԕ,}PZ�+m��Ǻ
�x-$�hj�� �PƟf�L��YjwY�r�h��c����;�Z�e:���g�d��E���Zz�Wn��C$�[E ; �u[��$M������e�S5T!*AB�~g>O#7��V��d���_�.�ȹ���<�m���`��o �����6�����2�*c�.��,a�y�B]ص_Y�F��3
����gu��	<�Lo�2�yu&�G�o�z���P[�W<w��9���M�}wH�uTa�!D(70������2q����]%�i�ll���<��
�p���|¾]�1�X�u�_���7o��|�R����.׏����R�;(��6Z��?���-&��!�hS���r#�h=66;F�05{?��:�P���(�KL1���X%��Y���`�j���s[���@�x*�-�^��2���s����yav��B%����x������R#�7�l<hg��tnyHlιV|܅V<z�m��U1������A�����Ze�!�L�s�)S�18=m:���Z\���^��+�}��Y����hH�>ˢy6��E�H���|�`�;�k�[/���P{r�ھ�=s������eu��Yu�7����|��"L��c	4N��uٹ�zḷ�A\$bT������H�L�	֩�m?:�{3ߍ����ax��I��hA��e�E�`�c1�9$���鏠ڼ|Xf�`�g`; �0�y����^���Y��_Zr��kFn�a�拘���ˆB���pCoDKe�l^l���+ߓ�,���2.��~B��x�I3����زe�d��:�k�{�t�6I4ㆽn6����Y�9���VU^�~\��L�O��>�`�!�>0�e�{�T!K�b�����v^/R��?�}�&��}F9M�:��ƭ-d8N�k.eºS!�u�W����RB��p�0���2�����w(f9Vbx�������!e��U��8�7���
ߜ�ä��kf�����vt���03��<~u>��r�I�����t��u��h���0A��(��o�Z��n���~#d�bo��� L+��>պ�%��F�,AQ����O�6����%Z���R�H�v�+T�b������yM[��$i�A�6��Pc�\	O�cD���jZ�����؇n�)Ga��D�a��.�邼�GMj����5�����/^���&l�7��M0�\�.wqs�m*����,(-%���b������Cr�j��P�p�5�4q"GG�������gM�0��y�*w�8��9 b)U�|��,単A�a�J+�G�춖�LX�xY���V��o2���������Z�|�v*���v?�:PGI��8�k�a���l��a�OmyY��?����|썢"Td/Ky�@���?Ϩ���S�]���2�X�]+1^O/h_���>H�� �n<�G���� ��'�0	��?)1��O�6�</W��w7��"����hCH
%;��U��TL3�P�2���Cp���9�P���dz8T��;q4џl̈������o�d��)j;O@����O5xL�x�T���u��p.|��������{�B�}�d�����ꧽ?kQ�o��kyx��vw�ӥ�*�:lB�U��Ѩ��|	4	��3�^,�s�#�H��3M��͗�8��֦�(@�{$��L���5LY�$�9��j�սhQa# ~��f^��@��߳��?�}�<f06�OzHsLz����Ķeg��Y�Hx�`_�'g��}�9�f�mߗ_�cQ�X��M2�#G�+�=+3��3&��v���y�h�9�2�����
b�� e �5ˤ��HC#d���HE��0�##*C�Q�ѷ��!�c>kS8\��/pd��o�#���r��?,��սh����7�i��6�y:�#�����1١d����ߞ�V<,{����n_�Nq���n�W~C*v�/��٘?�;��� W���0��{��)v�)D�ad[\*V�ǈ��Cx��Q��5;}ѳ�r�T�����,���_�9���y]�������A�zf.Jƍ$�LYb,ꆲ�L�j�X�i��/�4J�4�����z�Ѧ�݉'�_�W����ؾ#����npq��"�i�X��`UU�)e=�u4��J|y���;����l���Dɉ�H�?d�#�*���Q.+
X+!�ꥬ8r���������%m�H*��nhKӳCnA����)	eN����b}�3y�V���ɰ�"���!�֞�cj̄�By�w��A�m��l�57�\d����wK�\��w�-���ߖMFgѷ�Ὕͮ��%Ãx�o� �֓�}�e��x��;Oӝ���,�g,�$���S���_��r�K�3'���?G��_}�ok�z����
O�Z9��$��IDa-m�i۝-A���̬�����V�b���?.�<�cg��C�j�������m��h؆Wr���|��dI�{�����+i6n+�[	��0F��[+�<�s-$�iG�`-�qAm�]���&J��ȿ�>5b�@���6%:�̲�Q2��$�.��Pg�3Ќ�|�%X�m�'+|�m�w���u3�sʪE�Nн�/(��b�V,��%"=�b#�y��Da!�:ō��/�y�_h�D�6�\��3�cnJ�K��F��&�_��)+��F<��f��y��w����/X�_z,rYÈ��(ۃYk��V��(��>�r:�9�Ʉ������˺k�Rg��Ƞ��/u[7����ɓ�i�qڪ������K�pIV���:���h�u��;�W��:���%.J� ��\$����|���q�ъo�)�j����*:k�{�UP��F��eV�V�;O������@�~�j��u�?�+&j����/�2.�U����>e/�J4F'Hh������J/�ݔKrrP��_��M� ��W.�x(�XX�H�6*��A��.�B��
���^�ȓC���S�*��Ҳ�d>�Bǥ?yO7cC�d\��N�Wn-m�RuIϞ��H<����͐Oe䞚|0k��{ȼ��n�?��l��;��60���(�E��OtB�R�E���R�o��BBCaD4?��#���qg�����:P��_���jA0O�.���7<��d�1���@���v}}}�;hո�WX��^����xm՗�>w����l"�)�ܫ*��S�W�Z~�)��c�#��A���x����E����]���:n��̊D�+[���e�t����%�#����+�VO�H��7"�X���ġ�}����>���5�BB�u��t~/�k����e{O�����>�WȺ��8d�`Й�:Uͺ���ڇ ���-�?�J����L�gd���%�m�`ѥ�_J�J4��y�-Nʖ����#�u�{l���I3��jx"�9,�b���E�r0/V���`[W������� c�_{���f�ũf�L J� ��Ε�H0�,:��c1�@m�:"%d7���A��SgL���;���P�L���V��Z	l�k|����X���������T�
�M&��3��|��6�Vq�g k�P��s��ۙ���Ȁ!_?@5��Ϳ���@
�O�(��rbDw�j?�O��ex��B��e-�A��ALD�V5�[T������4=�Z��>o lD�;<�x�������7HW]H�^>Zѐ;��{e�Ϗ|�]��DC�=a�'T1:��#	:
���8�x~�9�]�����D ���4ڴS��&���ŏH@����-�
I>�įn�y���2�{4ɠ㵹�2[�R�{(�9����l7]�3�����z���?���������L�s�_U�Wxd�4�ql��;���ӱ���͂� ��zx��5N�1X?��kP��B;�N��h#�15��6A�k��zV0������Oqݰ�6L�e�At#7)�]�U�"Cօ��h�B	��_ޔ�W�r��'�����U��S,踻�P䵠��Hk�;�
���c>][1(ƻ�~_%�ZԄ��gnq$��y��9�$��J̖��F�#�����!���)ۓ)U�e��'C��c^�3��:|���]����2B�`��:�S�(��*z���ӻs��M�H�otm6 �K�8�)%���@�JFGw�	��p5�@�ǉ���Id)\6�
S2�������������I�
h㙞��K�7v�A*_*��t�ݩ�@`���*��ȦK�rp��p�I"�1+����?Xw>�3�Z�n�V�P1���gO��'~-�~����B�!n�K�Pb�k�ASkX��S}�s�j\���e��g�P��@���������m�� ��[��7�м��λ+�{�?,��� 삢��	(0�5Hiu�X�w�xK�s�GTc�'_�M��\\���u�7|�L܄#�t�0��Ӌ�>7�~�F��wr/3]2(�*a�n9�)�	�{w��L%�����L-,݂����%�%,��S�
�f����o>�7�>w
K���k�coMx��,8�"����k٦��4"�'���Z�?�}�sc@J��}�ӵ�޹�:v�T���C8;��DEᣱ7��Y� t�ĳ&��Z�,w:��;��)յLj=�Zo��f.y�.
��I;RCu�a���)���cA�u�ZD���]@��A��퓁l�u���R��~B�_s���i$�QfFo؏���_ME�I�>ˢ���GLA�NX�4jq?��c
#+����q�J��V�.,J�bX�"��y%���� �xT�7{kKB
2f���̅6��imIo��PO{q��ũ9<�	�Q�Ŵ �O��q�L;A�e�oh��%}��Z��pys��
��|��M�8k�Z��� ?+�_���k��|��÷Tg1�{YO��_�EwT�vr�BZ�(CA�T\����ne�RJ�����ΐ�#�]=�K�j.��m�n~�O����U���o��x�t���=
����K1W��ˎ�Hܬ����4)�U�����?㵯�J�)��%.F�:\�e��Tmq�L��/`�`�ձ,s_�_���	�6� �c�d���Y獢(VqSq���m�$���Ã��'�T�>��z-��'�&>`�X�}�b�ų�H�������w��	�]�
���:H;�nלQ/n?�l㾐��d��O�l�����-�'��H���`�2�&O����^�E@Y� ��!�?���%�v���c���a_cʼ�m�2?3@|Ց����	�{ֿ�0OEn�Py�����XLӼ����aUu]�(�����F��S����n����;	�i8�t����������1ǜk�������SD!߅�����#·mp�@rc'�����*�w�b��C��b��I����$\c�o�h2gN�%o՛ɰ�~��Lm+�r�<��b�/��؍s!~!憑���bg]{�8�ރ�|�m⽇�y~�ݳ�vʣ�S�O$�;��a%�Y�`0u����1��>b$��L8$H`�'0!�7v���Aէ��r\!Y�Z2�{��5�Jd;?U��4�bn%p0�4� �W�I#�F�Ӣ�(B���X�r��V�	'N��L�ע'�h�`��K���4�������kT�3Ű��x�����/<�����Hp�
,�FO,Sw��/���w�
?k�IV����BL����r���e�:A����;�K\�0�����a���?�*��<21� oxY����++^
���a�����6M�>uC��Dt���I#�A��&b�M68 2�J/���3jT���].E)�͉4o�cC���C"��`b���3d���k�%��\]O:���Y�5@=�Z�^py�����5p$�� �����Qy�?�z0f�7�����b�2�*XS_�p�e;K��H�b��"h��h��	
��f��x���,#A��ظ�q&���W6�?��[�P$oN����z��s���fl�<uTx��l?i�W��w���乭�X��GY���k���JR�)3����Q��S���uR���hQ$*3���؈(�d�>���lp�+	�,Tm��sK�CK���z�q�Q�ѝ&�|`.	������n�۴��#܆��dҞms�Q�Ѕ��X�8�n���M���}�u�1�:�~��6G<(<��B)H�3�5*(ksQqK�'����J-1@�t�;o��159�������-�����2���N	�S��$���}g��D�%�y�r��@���"->8���e�I%��@5�Wuq;4#~��	|����I��W!.��x����gW�E�����������ɸ0ZT��ONA?ǰ&1�h� Ѧ��uI��gHoG��V�ܚ�"��o��=�MRWIW0I�x��V��'�T�x>���Ä�{%"dN^��>J|�a�;����VԵ�:�i/����V�����y�z�V�<h��iƮa1_�~ɉ=R.�z���XQ9�k��͹�VX켓�w�������~`AL�*Q'�P������k1DH?��O��/]�H�8�kX["�=�;�����ͻaY,<x
�4�Fy4;�Zk�;�+!�r�� ��0'�p'���~|���/�������}�* ���1a5�*�ɦ��/�H��E�DQ��5g��\GuJ/�YwG��S�*N��٦�Pfէ0����t�(�Ǻ3�����BA�I��3e5��P�+;1����mND�BS� �I ę��|y��B����[�*��ɕ��p YJ�_Q��ۋ���?�+��w��^Tw�|bX���\��Hv�j��_�&�+*E(��m&�>[6I�$��]�(NnK$���D��C.�S�C���K)�X��Z��Z �I�W�(�bb�{ӏ:��zw0�Ҙ����YIOc��лW����c�8G��ۼ{����Dr��I���e0�y1����ԉ4h��fP<����I�O�} ��Ap	�}X��K�K��27Hz2���!�v��2	��.���$�Y�5�;es����Q�����,h{�7�*�A�q̷��ҙ�U��dT�p�:��$ÀֆLy��Ӎ�P�ͬȰk��%���a��?�fVɪ�Pe�,���%����3��l���<+�Ѳ!p�oh56�X��
�����i��G�OI%{*B�/�f�^�qd�w�EYj]^/��3����������)�i�%9�����ެ�b����=)V�f�m~���q\>��0v����Y���)~�I
�;6�����E&���ϐ,��W�4�/��y�̱�]��X�h�� ��Kc>%�R<`O�^���׌������1��w�*2�p/�-�RȂ��cͲy�z���AQ@�E_p8Ep���/{м'�T�Sӿ�~�hDPCbH���;g�?`�s{��Z���A�ѿb�RU=������J�O��i�� ��i���i��s#�=�������n+��J�b��EO� @c��髓��!Gs�04��Rj�GШ��wû�u����e��/+�& o��[Y��x��,�♛-����pvP�!?��2�QM�:B���Ârn3��|��B2�c��7� ��ݫ����p�n��^C����؋��G��y>͚NQ}S|����0�dTe��(6�L�?u��M��9���lE������Ӳ라��oE��!������ʢ����We�S)�p��GF/�+&̋�n�v�s֒����
�'#������1
T썑5��A�oGz��*B�*�>�K-�T0ڐS	
@_���$�S�ܶ��b-fr������i�+�/��� ���û��uH.�E�KP�"=s��`!�������
N8<Q�&��s�9����m��8��J��.��
�����j;
ze���gWU�<n���ִ0ە7��1A�Ր�#?+�}�l'�>�́�D¿x{�皛��ڗ�{+:"W���:��E�h���\�!n�||K_N|S!����� b�?���m(�]�~t��V�F\�IhJ��O����j�O�Q�[�0������=�[�EN���B
��U{�-���^�R#7�b�|J&��,��9ۘ����ͅ2=��4�ԯ�ԧ��gfB����ś�>d��0\#����{��A�ω����O>V*��K-\v���=�ш����Y���)=��?y!{ �Q!6&(����y<�CZ���'��y�hj"�Jl��A�&g���I��{���EU��=٧�ּ�\w���*/7M�Fϟt��΀8)����^���@�:�7�7�/1��h<�F�Pt:�b)i�1,����:�z�AE)�񺁅��%Q1��a|L2�D/�1�,j �Ԯ��� oY�Z�YHF6��E��R�ݜ]b c�\��G�����U�C����V��8,�)�1F
�s-J��5Iq�B��dUI�P��s�z����*�BAfoݧtj뗖��K'�����Zq�oIr�}K1�d�~�P��h1eIB��G���/	([��f~Ƭ�
� ���c��ɢ�
�����G����M��*��?N�۸�>�yr��ڑ\J=>_.�@��D�����$� �EUn5�:zE�0�p|A�'���PƜ��e%��'�G�E�<����sc^�ߋ�32���c�!��$bI�:���|����Y���ެ|�#�R(��B��J&m�yF�4W0
���;05���j�o`��p�ڪ��@�&��������t P8���QHd�Y���σNu]�b�j�����q`��O��oK�l�!�5�"t�G��e+�:����/��g��Z ��!@�ʑ|�(p.BOzZ��:����Gm�ɽ�J�sxM@����g�����ԓϐihI�2���p?�քK��7M�x ��ֻ�Ԡ�&�o�6��L�+Ƴ��P
��?-����$��gXv�E�-HP>����U�:��MJ�(}����WCV!n�Q�=X��6'<'��l�/*�[K�7�~	�ه�
?złP5Ӻ���f�}r:HKt��![���j���pO��I`M5�\ǋ7
�#_˲�r��n��ک��'�'up�>�����>��3|����#�o��D�Y���{� �k:�r��0�)���"�R����MU)��Jl��S��;��ioH�]?��KkW�r��}+�v�����ىT(ޅ�5�ʹ����"�Հ@R(��P hi���j[��#�7�0�c6�����\�hP���}1�J��sa�j@�eCz���x�Q�i����KNS��j�V�l��п��x ��[��I�/�	i��W�O$����~I���͊�O6࿂�k�j$��V�DãdJ �L���ý�yM�/Z�R[�Qٵ)gVQ�I���o4��88T��� �㫿!��>F�#7?S���4F+�#�<�M����ġ[�A��b�&@�@|�(��1��/3'�j���Z6����|��@�<�6�s�B�})Z�X��%�a���%���DR�!+�I��7b4�3�����az}��_@{.�s�ia�*�����qX������G��	 �&��/3� ����A��2AbW�s���-va,��c��N�׊&���;ai�^/'�Ǧ0��1d ��~)�#V�`���A���5���?d�[So6Kd�߁����^�'�9�&]w(o�%��xPL��RidF��u�)ѭE��l.�*�q�Mo�^G���Q�����
�Ь�{�ʀ�_�)�7����ķk��)���0U����
"u4�*�"���W��Nz�/eř��e�:�_6���ȩ,�ӎ\�~5�{$�����:�/�.�����[��f!uH������'{��Z��!�G<��
i�\?�P�v���> '�%��y�"�Ev������
� X�$lr?"��~�e�D��ȷ�"�k�_����,�uh#�>�N��@�������D-�z�Z��=�QQ�;���TzT��|�\�U$�G}��u?�[�L��0Ѽ�ǅI;Ev�TT�F�m3[B�v��Oe��e- 8J��=�D�~luԔ���Ǉ�I������}�ͽ:.)�Gm��?��I?(;���,}�	��}R�jY� 6��� bXb\�j�A������-ژ� ��O@�&��<�#8X[��Gz
��Eg>�n��V�\`��/<b+�E*6陆w�#|��o@��[t���M�*�0rc�5uV�����W:S��	���~��+��X��K�� F49�:�T|^_�[((�;�EI���p��H�����ݯv�J���!sh�N���%L'ʅ�h�\�\��/J�(r�מe�h}�EӨ)mX�Z��U�wU�&�o��P��
�`']�W=� .L���&׊�o'v3I�Y/7�!!��D�2h0�Ģ`�	�.k�R�Fґ������>=�������K��U�6cA���ׇ)|P7�e�3,�������ҤJDザ���\��-ՠwV~����P��Nu	/#IR�.� � 7R��$�����!��K���$.��X��Oa�X����Q��k�����<ilU�l������+�Z�!�EP�&�*,`*�Ͱ71�4oy7���Y<���-Ʊ+�6�j���b_,�E,G>8��Paa��S}���Z��B�7� J���Ux��MU��������>��� }M�V��D�ֿ9_{q_H����J$������d�S ]�Pa�l������
|x�Tp�=>[��ӭ3 rI{T�5����O4�s�P��:w��f!�a�8�A!v��}9���*j�{��խs��*�\��A�^V��TG����G�'/�􅘃ฏ�����12]H�=0]Ki~ǿ����z�/iK-�����Ađ\s����=��e�s�����z{�ˠ�>���b�w��������Fx��� ��&�
�N�'��a)\��Ϸ06�(����-6_࡝��j�?��@b�J�,ׁ?��r�AL��u�;@�t��/*O�R�p�Cw�!��4.�z�m�oH�W��ST�Fo�XMi���5N��l:�>♭�7I�
(�$�����> 6�/ M�W�x���o�R��8��9)��A�P�uY�5R��xeZc��N0��_�g�B�#ߩ��$5��\oR�M���X�]����8П������TRl^os�,BL�}�q��Ⱦ��T~"���᫠W�+��6����I���)�N� S�]�a�;��$���^��} �T�9ej�>b ^b��Z���v���|��$�}��ΣCc�Sm�#��~�Y�V��_f{�z�
����F0���}�:���i�ˏ�Oʱ�,������^��D����0��� �Ȳ/�|��:M���nn���v�P�M>a����\v�5_��6x<h�@;���PfI�-������l�^�=B�{{�6� ~���I�!5���:I,-����
�����kAД�J�(�x�JN��/�W�-+�A�ݽ$E��l`
F���	�\���9������o|n++����YK-��L;����E�]?����c+�_cYjb��/bG5ZY�%f�P�F�&|6|Q.���y�`��ȭ�C�wU�thxYS��Z�u���b������
����^ap��H��J��9���`H/p��獏G.:�헳
b�N|@y͡�@�~�X�z�֔ u�G�B#v�0��oz^�wR6��/�����v��t:��f,:X}|�r�w\���!|��� *3{gl)�z�!S��YH��W�ȶS�fPBg+v���"�!2���M�F'2�!0% ��Yuɯ�{���ݽO����b,oa���D��^�(�|��J��k�K���)^׃�OWQ'ӵ���̷�c�
�B���OE��旒���_����<Zɚ�D�v�evά�
���<�c�(�h��gYzĕ�2j`Sx��#�����U��������u0jD��.8�+�����l�u�+�@���{�k��[�G
������v�Ů��Ey��<P.Z$�B]��
����r���x[Zj^8a�������oe5���,yޖ/�`.e�ozH)k�'�+�B-&���1��=#�@�.��b��JT/ɰ5J�;��2��]�>�ca*� F�w��t�\(q�%U�.UYZ�U��2�n�Y����u$3}v���2]�SWQuJ����]a��*%�$�g��]��H�l8[��w�w��H]�i��Wi`<pf��~�	OYjl���������l+�a"�n\�^Y/6�}}C�}�H
w��lV(��ɗ_�6��M�sr[��~T�K����2�����D��R���_��D?�"`@ G���(�pɂ��ۼ5����-�x�꿨{�	�Dk��;��Ex��R�צ�Q�\�=�V6ʢ���|��P��gd�(R�x����u�����X�w��v^p��Y��>c��s�NG?��H��ʊm�p�YP�H��N|P@��o?9Į�ƸϨK�Ş� +�,�d�=4�n=P��L�dQ%~�}��|�I6z~gUu��p����z)Wo��I&Ŗ�Bs�W�⟑�GW���p>�ڙ�b��z��b9I��D�45�&JB�����h��2A�[`+3�@��B l�7���"Y_to�ϙ<s�$����b
r{=��[ȌѬ�4��9�ù�=8<�;�8M�ݲ��;�ؓ�ǹ�o��Gb��|����֏���C��������@�?�U��N\��]lE`����E]u��R�L�/*�T|�_1fG}�c��,u`|~���<o���ܬU$+�?[���zb��k��m��q:yݷ+��J6�!ȗ�3�
Ė���"Xj�y[ ��s������~������`&DP��ޛM���s����*N�퉗U-�X�]�P,��y}�����g�2�$�tqoV��ǿ,u�[fH�/��Nu2AZT�%tH���>y�J�ց�x���3�2���g���2E Ěpz{/'�:؇׬3���f=3aBG��Gzu�cC�����wg9��;m�-4�(i�����P.4���wѾaZ1���@�w��W��Qi�,�K��H�~՟Kc�!�iM��%��L��HX��p��fT��B�$;�h�!���\K0�{`�\�uۓ��l���J&������������N�J:Y��01��J�l;+�9l�Mx�:S���r^�PB�?(�D��
���R���!⾫��ܜ-�_e+�z��W_r��t'�Ih������q���Bڮ-� ������{�x:j��a^�E�(����MQ9���Rl��#��%�RlƄ��$�B&i�b��ߎ����]��3����>�WJ-��>�֛ܽ��s�����&�9dJ)�ة5˲�-,d`EUr�еC�����GQ{���?�T��%�g ���Ho��b��wn�+[l��2���Ҝ��ϗFp������8l��&�.,:�����!%ߙ�L��RC�<pa4��; gW럾Jn.���uWq�5�T���r�h�>�p�*��9%f&����|���M��XZr��jzB�['��B�c}�ň�j���.�j.�\+6,,bb���#g�7����z�	���7ci@˯B�:�`���B%�#����l,=&h��n�mCף��M��t�n�xh�� ��L���0�	��~>���F�W܊��Vf�T#)� �԰�b'wz��U
󇶯a}����^J�/�[$���������K$��|�l6�u3��w��.Kh�|4̵�� խ�4�����Vk����c19w��NdzJգ��3�2ת��q9�����>��	�V���OEo>Dƈ�!�������֜1J�a#����p�{�^��0��qr����0��p��,�łH�~����r�81q��n%^]�!j�v�v%f16(�V�{��D�k\n��r��*��n3�C��y�X�!�`�͵g:�>��B�a_6��К"%@�Eitم�n�e�u��������yb��F�K*�ԭN��p��� �"������۲�
|�+��ޢW�:_XC=��E��uj7�~�ח��J-f˚Q�j�H��k��z	�İ6���N(õ����4d#����q/$7P[3;��I�o��W��Hj�#QOS��`�N�\k��J̀�_������߅�%���,IM��dHd��@���C�M|�ˀ}�WS�;�|^���`�U���g�|�/���mw;�+$n͎#8'�x�f�0&���1B;c��Q/���R��M�KǴ]��]���o�:`�f��A䷠���.�������g���f}y:U��t����m�Mq������Q��,�g�E����eƈP'��Z���H�`'�C�c����7s�%���4�VzX1[�`ڋ�cI��#�L�$��t5&~u��'��%O�~�g,m���x���b2���]��3,�d�Y5[her��]�ƄZ�A�����w%�����\̝Tև����_4)���4�7��!$y���1�:հ�����e8y̵�y���Դc�{خOS�l��m��@�Z�qHY/P!�s/�10���R-j5��	sLx1�?���e�C���K�B\`��܃~���K}���^C�9���]�)�t���1�j*�$�IlBɡ��!��y���L��qc��I�a��~�>��6H��L���`m���Z9�?2�x���i��w����5��i��ĵ�v�l�a�>��3�EW����>�}l�v��j�*���C�V�
�;���ٰ墼 (�cm61�H���㘙g��*�<��y2q�O�aŒG������`�RY���i{m��}�y�Ș��x��O�+��g��SJ=w��'��(|M^��*�H�.���wK>�!]�t��lϬq�81�������Z��D��&+��*�^C��N���U3r�H���w�4�ڼo�#'�����Z�M9.�m����f
�)m6'et��GL5&�k��,�T�^w�S���4�N���N���!|�2F�=�xܗ�8(6%t��V��N C���Ah�� u9���~��y�C�4n�������v�c�٣��MG���oG��`Kߙ�P�YgH�|���W��W��ƀv��^tækq1��Sjn���5dp�敶�͙.���w(��"�ίF}I��Z��T��h(^K�E2=qX��'畞�\R�	� l���Sz(�n���a�,3i&yc�/gg�����H��� J�л���՜��-��QC�)^���yuoo=ws�5zB8y�s�ī����*�#l���Ͽn�1o����<�#�f�$�Q�HXg\��1��9>��g���\]���h�9j�j��1���"�|Ox
�^�N`�S�t]�F �C�_�c�d���o�\���W}��AÙB&t�]�*iq4����:���>���?����#W��k�Z�`�V�.̯�*�]
L�a�mM�-�k��NB����i)��e����U5�~;,��;̯�J�U�quUD��:���
ϣ|[���}��ɠ؂H gy��\*�LH>KL'Jj��"06�t�-+Q[����NQ���Ws�n>^FȎ�]�P���d_ȸ��gm�o"�HX�7�g�wg���q��}>[���p�:_V/4��f������6	�ġ��Be^Odp���s�W6����2�%���$��Nm������-�*�ԲN�Qp�����'	o�9��aR�����/*b��V�2�.��%k���y��$+^�r�݃�6�c��r��R�}����9���$f�d�]ʻ2�����і��,-e[����ɼS��Pfѻ��-�;��o���k���O��C�+x�j�ω�[���J6�W���t�{�͍���(���!�_#��SkJ�E�_t�Yh'��>�D_i�����5��M���@�8������_eO�m�H@��od��=����RԎ�+,�r���g���@�wJ���U�`�/z������=�{���4;n�����WN|��J��*a�_�ƒ���n���� fR�Z����Y��}���ߜ*#N=�^���:�Be�w�(�9��� J��,��Z��Y8J��<�\W�\xh�p��,��.=�&6�L4<�7����
j`ɬ�ݍ���b�lf����F�q�Md>�����0�
����7�֖��0�֕C�����$'3��f*��Ӷd�u��⋑E�3�e��X����&�z���I}���[�5>�Si���!�
1�r�UDC �! ��O�;���b�[��rڑ��Ά����#۸P� ���c[� ,�x���Ē�Y�/�^�`���Z8�c��_]!W�;�0 M{�~׉��4Ο�Q4�Qf3u6�k�����	. ���8ٽ��jOu`;r8YE��D��Z:1zU{�	S�a&G0�����AX���s�ʺ4��(K+��Iǡ��u���;��m���;G����qd���V��0���3�a)��]@���b�	K�p��5�ٝ�I�.���-��ҷ\-,�8��D�R�Q7�����q0��s��r):�L]\L��vey���DFG�N�Vv]uZ�߱��$�^	����^G���z�a驠tV/��a�/����q�������1 �1�2�6�=/>�m>�O�z"��%�f�7k�H]�oB^��0Q2Ƹ)�7�,Q��X��G]c=Z_�7h��$E7���#��$8#�x�~�:�8�3R~���M�>��ӈr�K�8V�����6:m�p-r̘>_s����{�e�@��h�����>a�8���MF�u��/&	�������dR���G��a;I�ل�V��춣��n9�+N��"ˑ	E��g���>}sR�����u��k��M��#��:u��axƂxt�_�-�dp����w]��uH�S�^u�+�@�:���(�vwʬ�E��c�~��V9%iy��:CAe�*���:Aam�agq�&�/J٦F2V��"��2��l��ڳx�/W����H�w��n����W���3����hr����j|�j�_xlz?!f�@�D��h�2p�\;V�G2�
}B�a�Ӽ�\�2���N<OITs�"�FU�L���yq��a�:���VO��a�ol��vJ)Z��e��`i�����Ze�{h{/1^�����F�Ϧ�Z�S���kH�A�)���B[15u���S�;ݞ�*~[(m1��-F0]� �i<���>p����Ԍ~�&��?�����]�x�Tt|8n�eZΒP���h�;��Q����8�&��wEM��`#1t-S�e�)�9���{�����
_�gI�̰���cx��K�1���]D<U�XS|�/�ғ)�%/�q��&��@�,�?��w�E�I��͙t��XL�����V��沒l�s	���P��α�������3���nS��\cq�|�m�������dZ�ǭ.����r�j��rkY{-ɜ�r�Z�,N�L	��� �Q�E�A���HFVieX�M��9�^F�M��U���D��2駪C�;���{T��ϔ&My��Qޥ��\�74k���h�}Zqay�?��;���T7��qz�ׅә;�����
�'Xn'[Rj�z~���,�l\gsãaK����	%�z��t1���I�C0y��.jϸ8�
"���M-R�ù���U��#����yg�I��s_�_x���Y��|�pF�CKk�S]�� ���i��(�J��W� ��aXb��z������s�|f=��)^���,��*��Ɗ��ڵ���!F8ʴtb����C�-��\��H]��~���@��A��č>�i;?Ō|c�\\��CbM��������EZ]2�֧����>;\�h쌗�ґ���e�<��������u�_�~H�8��Y�^l�I���j���D�^(3#g���(��/y�nscHl�J+��Oy0P��/�ˍ�θ�Ԥ���:'>Fx.#|&< n/�����9��aV�X��X�?i�H�*�m�!���»,3�1P!(�Zq$�p҆�0����n�)�^�-����[����CJ�IrT� ʳ����r-�U��CCT��0�Eq���Y�ow� .]A5k�|���>xC�׎UX�$Ԝ�Ր�b����"q�3�� �,���k8�w�-E�Ϲ���&����j�	|��v�H��� F�/��9k�'T5:��K�f��ēb��F���=.�Ն&���:�Os��u��AG	��Ɏ�۱�L4_��&İ���f.[Pj��6 �T=pXI�E�'�,g屫�V��vL*/N�D:���Y�1Y�g�8�����7І��[b���#J�a����l��$�oX��
�(��<d>g ����׉�� K�U,-��{�r�Ey�!z�A����,p���ǹ*��w��$?س����y����b����X��-���L��=b��Z�q�yx�w���B��U��&�߮�
Q�[�J�f���?�j�q;��qzw��9�\�a�����,�Ot!X
T���Z���� "2�ea'�Z;�3O���ϹB�}���Qh��u�1�c�<��f`1���9Cv���[���w��<zKo�"����ԧ�ex�i�ɹ��y˥Hh3+��8䷣��'�B�?y������pT��W	}�Ņ��beq�N��M�%��b;��� �� J�UDr�!&��GD�>Fd�JW�M��d��_��o6Ȭk5t[a�[~M�h��
�6}qDc���I�����/���Up�10�z3��&�o
v���+����-����� \�>D���p!9?���-vX̡u�� �SIp��������ٰ�5m��E�a��e����c��П��CVJ�b[.W�<���vϑߨ�Xv�{j8��,ֵ����N0��l㔶%�xM��;M��i���*�r۽w����m_Mf��c�l�%�+z���pa���M��w��Lo̿L-s_�{{⃿�����w5m����V������cП<u�UiÆ���>�iQ��
���g$MQ�X\$�R߹��BV��=*h	���<y�����c�k�_X�]���&@0������)�����;c1=�3��@�]�eg�Pxe�������ӟ���
|:����;�qN<���"Z�=��1������W�$m�I)�1���H�O P�|�jY����08�~:$i�I��<F7GOp�k����SĄ��6[� Y��Q�A��Y��`��K�����A*���W\c-�Ӥ��ӹ�У�`��˛�k�ͧTsU�NYz�\8Og�v$|ל�'4;��<)N����H09D���j
�8�eԵDG!��}�=��7�e���<sK6G�0�qbM��U�4��w�V�յg�A]�\��?����Ǿ�؟ $q��D��`��-���zcl�i�HN����.x�T�QC��+�qi�dތ֚�W#cb^����cBg�u@�P�w��հ�:��KQ7����sw����2�������Y}�E��`�o���zv�`�Cc����m��Q�۬8NQ���c5e������I�0-.�dV���xp*�h��p��I�Z���-�BfT%�_��8��R��{F]��k�������e< :�+�8*P�=f�J̋�����ƴ ����<j.ο6?���"��l���Y��l�}T��_�)m�>g��,��G�h��5I�5�sx��0���N����F����Z%,���J�cp[��)��RWT!�x�*|��K	/_� a��j�W_��C�dB�V�w�z�ֹ�	�S7�m�>�������FKZ�C�%�az^w���Q��2�̣����k^a���]B$��b�z�m[�4J/��^~ʈ���XI:7�v��C���5��6L�S��*Nc(��U�� �(+@$b�s{u(G6��׫s]9���q���Hs�G����O{󪫹�����hɢ+OZ�e}Ø]��Y�+�>r�9�w�0�N��AyN!q�MD%k�έ�F��O~L�u��h�d�b��]���1�X��Ӂ���t���p�%'L�7���8X�v�J�Eશd�sK�g*�ȩ�y�vd�>��zn��j���Io��zb �0�ۻ�R����l|��臠S�;8�N�2�}�#g��ѷ���5%�����#���À�m���Op�\��*4�7%2���ҡT(�|$�����I\{�$�i��׼Pώ�|��-d���_�r�����
D�W�OB��z���k�7���<�qL3�(��}`+ �+�&�������X���94���G}D/�h�j'o��{���w`5�z������di���"(.]yN]�l0ϗ!rJ���%�xH�O�t�9.��\Dkws�_��}�?�XXS��4���I�b#+Th}M�[�	���N���t�A��7΍�c[�9����i����K霼oh�*�j޲�\]"�aG"��"E�cr��L���b+K+�00E8v� ����!d��g�;f�ɆxK�?�(^]��;:���?�����6�5[r}1�a��h�YK�;n2GA[�ڤ�(���5�Pb�oq��s8�I�&˼��C*Z���_�8�JuC��<Lu:	��O8Cʔ����¸eX��ٜ�,������׬l$�B@��VA�u#�f������uX�_��\�~"��ߌ3*�z~v�<�Oȩ�.+��j�1d��12:�>�5]//�������O�l��h������Sⳙ E��r����֯H���[�r��Ǐ ������`"�������>>�Eچ9�D
+�5ܦ�I��J�ًi��j
�?U��!��ҕ{�Ѿ/-���eؠ1q�M�������Ӧ92SP��4ױ�=4n�T��ē�=�iE�J��ƺ�	��G�	�� ,+��77f�h��W��$&;ЉϡQs�f��\x#��p�O���0�������':*BFDA�(�N�M���BOX�pc���D;��yG4iR_Bw5]��z�2��J� Nm$j�
֑�x'�ţ��;����hc����Hڍ�]p�!y��h�S� �^f��\��͘z�;�s�tn9&����3yN�ҫԯ�\i�0�����C�ˍ=b�0nf���b�� �ax��� M��&�{��0�����鵐���G\��M�� ��}�A���E��UO��Z1����7cl�nO�`f�H6����k��Z��[�l5��&}F�
m>��>*�|�z3��n�'�YӜj���Ʒ�Н]kz�\Q��|x+,]��*�F8�����>F)i��:�s��b{ڛ�c@��b��u]�0�d\��g#/"P�4P&��`9���C�_t�Kdl$c�'7���"��3V%Y�r�����eG���}��֪v��Gԕ�����-ֲc���Z��U�aEn@�
-hQ9������	�;<��3c�f}��0�L����9Vr��Hi�wKuYܲ��k��؁ �F�9���k�Yn|�Ϫq��?�M���8x2l�Sy��a+��t�L�F����]��o�X�k�̐��!��jx�X�;�I��v����x�1�����k�#�d"�^J�7��*/�S{��	����&�a�pڋUқ��n�+q$�QG���(�H?eͣ���P/�Ru˾��������'�:(�vd�܂C$���?O	��������ak�$U��t2�ED2�A<��P1^� Q����֢^��!z�Y 0���`G��,��y���n(�JL,Py��m��|$�'�ՙ��c�8b./�j� ��s���.�巗���ǫ�L@��@&�O�<��h�5 ���NMd�E�� ie��~��Jw�.�I`[��,�M0�	����MW?2W��W��4��Ľ���ݵ�����+">�����g��*�4�<)�/�4��qP8�6�'��Tq!4F��
��U�Ɠ%|��!Rn�(��(�)�9���A�K��F�w�oN����qě�6��5B[
��9K���]�qH����
L˗����w&!��C�Ct��	f�EB��N�=Yd[b2Fy^�S��yު��G"��Ȏ����9aW(#�y��A�J��;�f�B��k��ڞ3��.j���e=XӋlIÈ7�f��5�|�]v
.]��G�WF���B��N!8�`�������������݃��vp�7��޷���Z�>=�U��vu�L����~��Z�JdXv'vi�a�]v�¶z�<����ɫ�(�$�P:���@���if:��ҙ�0��)]+�H���԰wF�����q`�]Wr���4{X��6� �z$�~��j�4�S�5�(B�Z��Z¯�r�ގX|�+-��"�j׳
 Pn���ϧ�5e�b4���.6�O��@��pw���F�{��{f����1��u�	��Eh�OWD�S���³�)����.=�0��~
,�(���P^�󂎰;5Խ�)	/Vc�>�������,`:����P�\2)p�F�~�u��z����
t����,'!���͵�Z����C��$�$��Q"�������h���\�tYًEz3^)�@aϥ��"�ԚmZ�I����ōz=��cg����"K/r%:A�5�p�w�M���1q+g� {�bҍ@8ԹO0%�fڙ���A�8W�p�g�)ƛ��j���'�_�EKE�Wi�A�K��"f*�{CA�\�wr 
�r��C��Le�M;M�?��Dߴ�Z=��{x[<�깳h�_J��z>����w�j�N#�����Wԫ���~�c�Mcz�ꪍ�-� r�Q[��g�5��*�v��'۱Z�� eDr�57�O���V�/K��:RK�O�V�7�W��!Z�
�OI��Z6�OU޷uK+������M�a[XЪ���vS, �;4�����Hm�pr�q]iS�y�M�����7�����A)���L9�ob����4��簄#���X?�n�\#��˯N��\VվF^T�!��77�?'k�LE���QA�p�,y��)���턄%�wXo�O�f���DP���"CcZ���0ts�Vr���}i�e��L7�C����w#<=��#�y=<A-
qOw�:�U�|c$��}�6t*:a���A��l�2��ی(����+�ց���3��Ӳ� $\��EQ�(g�*��+&]ƨB+:�f��z�
�xzV��A��<���2�/JG&���ٌD�<��M�&���2�"�ߊ��4�(O�)C�n�
a������#Y��	�A�Z��� +�Lk0��y� ��|Hn�N��^|������FE�(��T=��^���ằ��G �B���}��s[��^D����ݛ=��a�c1�5D�ޝ��uU����c�5��S����X͋��Ó ^�i��6,�%�W��o�ڽ
-�|G�C���H#��Ʌ���H�+��g�`����Ƹ�7�y�6���j&�}�P~8����aE�/���|3����6�$��bW��,�'t�!@�jb�qU�w��{ǹ N��b3"�/�K��㮷�υ�f��O^2�`��H�E�<GX��znѤ��v|s��d3��N!v�HH��2�͟s��p�2�a�����o�tb��	�\�t`�K�s�A���9riWu��Z�*�B�O�:`as������Zk��!��i�>��Lg�� +���[
�a1��
�7�ِ�haQE���H�p�S|��S:h�Y��_ y���C�o��Y:��+�1,��((�g������p�";䓃�G-7��t����;2�3�9�3MM�S7������}(�I�rV\\���$���j�_ތ��z�;q[�
�������n�95L�T�G��fd)�j^���&��B����DΗp=�x��>���N���q��<Ͽe��ͥ��މ��"�N� D�\�K7G���9���$���&�_�	 <��]�ş�����/ʓU���@��/]~sρ9��>�yA�lv�v]lB�<�;[����L�<���f,��d���X��wa$G%Lfٱҏ���(R��.A6�V�{��B�ǪA��ښe��@�Ͳ6m���?䴫��7�PR),.k���`i'l�ѯI&�G���S0�\xV�L�}�����@�]n�5�֊��d�������m.�[��?���������Cv]閠�:r��0�����[�b��<��U�H�*1�`�\�7��ZzvW�2�0.uHi�� g�vm���[��7�<��.��끢~Ø%Mg���D��\��y��p7��3�OY�K�a�.Mȟ�t<���Cq�.��/�+N׈�77}��?�1���Tp]��*!�F����Q�y� A��G[��Ub��Ɵgs���a�h�q��h�X�`7ۨ��{�]T�I�\��!F���H���H��E�z�:r�[*��i*C��vtFyz��#ukc?���>�ɗi��_�;��#�IF��B�4͇��fw��|׎�
�B�#��]�	�g�E�f���!"y2{��|�������@ �Pf7�������]�nb��0�s��_��=�*�m�W^��L�n��v���A��8/��ȷ� E�0��;��-��	����M��q�ժ�c~�9�����b+�!G$������ 5ryʧʪl���wE�3$�y=���ԉ�a^ĳ����/ՙO��Kr��z|���W��I�@9��k� (�̖Ki�T�2�}��hC�W�R�����t��N�����
��@4�vo��t��3}"����Je�Ϊ�Tи64��P���'٪G��߫�YY��>nWB�hٍ;�U�>��� �'f�F�Xc4��6C�g�Ӷj,�1�X@�e�n��q ���D�eOr��mG.��Ì�/����g>������#��L���a	�8\���T�&�<�	�׶Q��yC��c�}�ס���1����;U���S�~��*�<|�U|��գ���P�K���㮒��9w�΋Ȋ+�_*k�IK���+���꽘�Z.ܐ�������;��N�R�?��R��y��hA�\����=5�ރ��[?x�]T�0�Y��#�[�93��a����/S�@b6n��.*�<PǴ���*��kX/}��jM�C�m�����q+<���]@AG ��Ҕ����|uiʟ�Z�v��˴c�}��㗸���I�����ZY��}�H��-Г֞4ەZ��-$��8Ek�z��I���EBq������c��
Z�Y�h²�V�O'�/�(#�P��g�f!��&J��K�6�q_1�y���!�'�¤qze����3P��(̽�`g�ۭuD}����g-tZ�Fl$u��.�`�co�󾍺�F]�7��kئm'��am9y�#�r<c�*�������'�Y���I�3
?�Y�R��x	����^�����g[�-z4u0����<p�F���L�3r��ڲi��|���u�!�m�[��p&o����$�%a,��hi5qᭈ�%�r=�0���'
���=Y�-���B���qߋ=Ms����s;�:���16���l���/DAl��@ô�:(�@mV���,�u������T��B7�(~��:TW���r�;�Y�R&m��z��}kŷ��Ø�w:�c�������eQyh�A{�lV�h&?_�z} ���7�]\x�J�{S�M�#b�-XÌ���W��;|�� ��AN�����`Y������/N�y_>�a{�e�;yq���Oz���QX�i�{��ƥ�ꓞsrMUmť��D�qz���o��m��|�D��"��+J��(�/�V�F1.SF�U�$� �m���.�Ưb���~��WR^߸��qQ�p\P��I�����{���,)�7Ϳж�\��ݞp�e��U���^a@gf�δ+��Le�����:va��l(?�$	� ֆ�fHk�l�nl�v�e��\��k�y.a��I��4�gY����tC��kҢU�eh�ǆ��[;��{~�<cW^�e����L�Mc�Y��#}ՅUr��f�Tߩ%&��������T���@������p����WDnc�P@PV�Ҳu��m�}l�-��Q���ޅA	v�O�4� g�@�<b({-C}N]� O~qV���c�!������ɅB�U��������C	l��#�32,��g��c���#�!�4�$� �F�(Z��yHY�@�Dr�kC�T�
*+s��:��S�����!g5��R���t?Ժ�.�D!�Bx��I����o:���\wD�EB��mߎeFvV�s=���B��/2��P}����D.��Gl�ۣuk��p�"����3G5H����op]�SY
k����;43���q��(O8n���t�r��5�Wswb��ZA��[�Q*v*5f���"�x�G�j���E��K^
���h�4�+u۶>q#��^y��z�T%�v"�k��@�{h�q�Jʹr2�J���/#
�GZv�^��B�K��p�}�AK�0/[=w-���"+���R<��d�-O�_|A����-�z�%,�=<�8�ȮU���"]�������Q��U�nq�A}����Ƹ���]�����0쨷%�A���e�;�^�d���j���,s۱�9��TG��mZ���8iDc�� ���:<՛�>���YGmr��h��_���
n��2�>M��y�~�������}��|���?�8���, �����y[w��)=�����͵[�t�a�}��2_{�o��6 �<�#�j�eh�D�\?h��m42m���ݚ�8��������iNV���F]ʹ6|��u�Kj}t߸U�i�q�Y�T]?掾�d:iX��F~��^�LBn4d��8�N�^�l;��,����9��lYz�r����ɏ�߽��q�XG.m��&K��*�e���E��|�?(�s�W�b����`a�K(��-����{��x���
#�+B���_u7�،����؅a\\�$��"�ۦ�±e-�ʺ���RkP�y"��d����u���lB�_���	B����q�H���<��O����M��%��4G�N{�6]����wEUК$�2ewhY�sB6�������[0�X yL�,#;s!]���N�B�v\��b�>����H�$Sx;����ؔ�f�o��)����b��>
��bC�8��n�
�
�"�5����uW�J�I�\�߿�>掘�AmG	pa5͵S
"�DR�%_��gI¿j��0{N�Y}~�Ы��x7���w]�I�/��o��\[tfØ���0�l���]�7y��W�x��-���6�DM;���B KL�����Z�^_�x�O�$׌�|����!�sG��`I����7�V��K�@����e�j����g|�p�3v��QAK��$�ߩ�S��]�:���.�R4�O^jOj:=z�d�`ﴪ�԰vvu&d�i;��o���՟D��Z޹�{xF��Za��}w����{��a��Ϩ2B:���ۯ,4C��k�l_�ZRBEOd�x��3<��P�8`��V{{JwY��{�I<C8����Ƥ>Qx��1����2�W�?_>���M�թ�~�7�e���yy���ܜ�m�����Yu�n}���3e�x�/�c�QY-��(�f���"�l���ͫ"L�n�^�?��"x^α��Mٺ�K
ҎN��Ę��9q��S��*-ui���m�~�[<���#�L\�<��� ���y�E:5���%�QN9��x���lA|V�)�GX`��N�7��<����AY���1���#Ȕg+A��ʟ�?�x7{]�P�K��j9�pY��O����i^�݋5}H~W�� ��-�h�<��o���/?M��[�f#�5s�D �ۧ�v��B仌8ά>����2:�j{��0�Г��a'����"(�Tgp��W� :�-���D����-Wp��Sg@��K �\\*!�
�2.@v6?K.5��ז~�+�K ,���mxub�Ϟ�;�y1
?R�u0�ܻ��Z�,���ڥ�zͺ��P�F..�zx��i��x�R��ê����9$g��Yjی�=�����v1u��#�����#��Z�����J�w5۝�=P	��=�B��e�?�$��vֽV�i�K-���G�$�p}�h�Sq�{��Zh��GI��*�0��#��#Kq�����~C3�C�A�(n�[&�(������3�)��_�G��<Oc�i\^����x-Y�sB�S�����Z�ɰ�4W�C>M�f����R������+���շB���@��V��H!hܺ!�����W�o�k}>8��-�;]mٷ��=�y[8[�r-�����,֚n��O#	� ��h{�p�f�?ܿ}����z©>����`"8��6�K؁�G�Ϋ!�9227���ݚ��2G���zͺW�=��[/񮗌�U�d|;Y,+5�%�`�Y>�������RD$+�S4s[�@���J��b�s'�\s�,�M>���µ�l��v�-6;��E�o*����z!�L@%*DW��G��hY�|1"n���Ȃ�i�W ��D���w�"̩�@M��,�.m�O���$+�D,Orx�Xwry�w��,�����5H�H��r��Fx���+a?�Z;�l���/((я�Ec���z�U,�;Z��xz<�(�ڶ�u�6��}���%�r�	��'�kx�օ6�4�.����4"0���K�^�7�:�V�` q����_w��÷�+0�w�ni"���-1_�ȕ��q��;#K{[mfa��:�}�7��э�M�V;v�<7���ڊiw|M�����~��Y������u�;�QKT.��k�����?^]�S�
bC��_fv�)�:of���t�O���</;�������>����/9m���.)��9{s�y�=I #WD׺>���t��a���  �д!��Ч�)_)�aB��~_Fj̴�ڊ����1��S3������kc;VKE8������l2ԗ���^kC�Hj�˕e\p�'}~*���fk��#w<��)k�^�:�~��鍘��?|�jz��+(���^�� {�6��4�|����'֛�Xo�UVq�WjGcW�g`*���_F��\�E��M��@��m��"l��3������]ܥq<��>TW�[���6���A �m&�����^n>��Ƨw��,}��Z����G�����FA��7*�Ɋ�f�
�>|Z� ��v���߹����IR�7T(����������ε��(2�y)���2�w��XO���hC71�4�7�%hƸ,�=�J�iƘ��ԩ/7�~=�|lp;S�qbВ��s,�]��{�qOY	��/C&#g��/��B�O�:���4���:Iu�?3]��{�^��\0_����J���$��OxR@�]-=����C�Z3:.�Ʒyu8�ʋ�Z��U�!�gF(.����/�͟�����ꢜc�c�M����p�Aa����P�̜Z�N���-�0;ut[��N�^#��zˡF�Vd޹plT�٣�S�i�������ְԀ�
�Q��U;������C��)ۉ�_42{ķ>�.�qK'����R�!�3Qh�/1E0E�߀��z��7N����TT�͜+�m�Ֆc���D�=�k^ZXkj6���������<���2�����p��Jh?aʨ>0�^	�UǤ�$��\��Cz 4��b���~�v�&Zw�<�������&�}����ڶ@��|T��pZ���TS�C�����~Ð��_&l�0׉�p|ݎ�P£�>�uX���񻥚7��q��I����:� i�� ��2Z$☒h���.�(7?[b3��^3�+sNñ�K[��w�nVѩA��u��&���L�*���= F���)h�)FG���ڕ�5aMKl�E���B���������j'�Ik�α5qu+B�~D�3ˣ?�����V��:���˟���V��6��P�x47�j+��lܒ�ڑ�9������{���峴F���H���m�F��Ow��ވ���emM��C�3#�z*�]��'mō���C�@�7�grs|z��k\�0��ἤ��_9�,�5?��g	���5�O1[}���=�ް�Co�FJ�1�� �ǥ�ʪ�C	gVA��̣b��'�zO���֙�^�*Pp�����a�i�qҤ�ѻ�f6/��2#$#�1Q]x�UC�E�"MB$t�MUB�9C��	N#Sؗ�)a#~IT��C�����] �'E�bf9�Į�B;��[��h�	�,J�ЋP��V�ȐV7�����l�=�$���$���*s�gwN��
�$�[q�C;<~�t8��K��0xk>�s�O�c0���b}�sZ)���R����.�v����"]�q�:��ƫ�~/J�\S�����S٫'�j�A'x�8��u؞�>�b
�j ��ZՙY伆|e�:�P��~\�וb�4�������tn��LԳ�9�A�VM�B�<�5�</�eLᙵ���g�@����}9�*�23&���Z�|���;�2� +)(���+���%�{RX��/c<]�t'�d�E?*�ڴ��g�Ca;D �?L��
Y��>Ex��!�t>6�_��h<���J�~ �c?�#{H��ϧ%��`�c�/z�ZZ����q��qk|�\��Y�� 1$>��!d�������8YN��ݕ�/�c��]H��?��Vj�uø�}�mg�r��Tɻb�|�r�i���µ�ֹ=6m-k�
�ћx�m  ��UF�dO���Ip�ZD ���L�o�/�zW�a�nւ	�~@��+ph�@������6ށ���-��u��L�~���aD��0Ey2}���ߎ*�4ǈ�ٕ*^a��N�K�����#�&���de�j�� 9C��^}���^~Qb���! �o\a�ݯ��~r6�U1DC>�f�)%����$��ǘY/����v��s�7po��W��3���v��j93��`��aR��Vx��D��='�䎛XyD���'�!]� E�M����2W�tխ��5��^�{(��4Uph�Ѽz70=���E'�{�4���=��u�;0������� b�D[�Y�(��� �6��W���	�ј�/֡��������m�5-W��G����&XG'{�����S��:�����S���/Qhc��I���8
��k��p����E7FE�v2*�a����X&�O��ZnI�~��kM��0�[T��.���Y\��{���@*�;wCCW���X-WUI̺M���{�'_I6�2k��Go����}L+��;FxJ�|�K��cL�Q�FĐ��f�ֽ��Hb���L����,2#!
+�@#-��Z0!�*n:k���^�ߠj�K���-5FeQ������q�U��p{�V�Lo.l/	9���̯��1�a%��l�9:o����.ͻ��̽0��K��AML�-��2JVq�s��&�
�]?ZX^����V��2gmv��79�xQ����P���PV=��{I\�+n�D�)g٤�����G�9�A�O �k����Ǉ���/@���*��(�g�����Ǔ{b��=��moұߞ��X?r	��VWꣃ�xy�6�9�s���B����\��J��d�[����b(\�V�]g8G����9?���6Ti	�9�6w�_^v�|�^�(j	�ۤ�y+��O��ቱۚ�jV��	v�D�-���լ�b}N��C�hbyS�1����?Nz�t=��!��R�93�\�����[IݻS�|�g;��]WwE�'ibj��h���2��R�Oo���z�4N�vO�)߄�J��\~d+v;�p��}	�įwT�N��.@�T��#*��yC�
��Q@6�ٶ)�-I��*<nf��J���rV��$I�8J�0��>�
{6e^�&kw��ӛ�^�ǐ�q�J�T>�m��!$ү?%��m2}SĔ�9v�(r�܇+�B~P�k!'c` �T2d��*BR���e�˘�[n��/?���]��&�(�PV?<��:�����#����Z>>
�yiE�\3�������8-UAcE�.�G�hH���1�r<ǽ)D��:�#P'���^XR�_qxˢ�:����[��y��A�-F�-�-Q8��Fء/	*��mX�Lo�E���L���D^N>��M��U���-�8��i��=]��J�K3�/�{[�5�B�%vW$�=
���"�K�_��w����7W ���Զ��N(���E���L �I����f�������>Z��Q F��!��I+�q|�~�����' ;�<c%pNwը�1�>ቨ>v�H�(5��x3#���ĈP[�����PDo�\�v#Ƴv�D�y�/�8-;"������:�~̲��D~�}*����O�'ei�pY��@�4(���w�v+σ�u�*��s���� ��%ݝE��R6Z�CzV�?I�*r⬥!1d�-;�Z��xd��;4{�Q�N�v
�z O�W�1�V���N�?/R�)���U��G�u�N�Z��TL� �qcc�q�'��ʁ��ɉ�h�~��ʀ�=��"�|�T!�zp%k�&�ʇC�Ɂ1<��bd>��"D��C�SQ\�@H���,A�X����nV���Q,����Tq�@s �������b3�%?LR���h�&�B����i;��}K�邊yןE���t��;;m��a�^amH���Pr(,޷��C���I����o�0y������k�i#e�Υڍ'�DY��_�������X�,i~�ɩX�W�j3���d\�D�]����&s��J,	�y�A��qDԐh~	"G<���
�ݾ��a���k��z#���7ǮU����oP^4҅�g{���͙\���[/�ޗ��E����8ݪZ#�M
�0~2�96J0�^������n]�%lV�ѷ$3���?�L��1�d�3��*��:!��[�ǐ^i���+��`f�w�L�b��⁼��T�B�\�^nT��	�O(��7V��]��
f�/!��O4YS�9��]:�������^����&]�:�〡��,�z#�]@1E��9h�yv�)�`��m]�L7�k�O�<�/.^�#f�#Q����7�PH\����y�В��<,�(�_l�8�Eه�Y��ҁ@J�zaX�O�c�5щ�I��J�C
t�g�@#���K�Fy��0�Nn�Cm�>��y\���[;����ľ*����Ւ]�9���U���R�����b;x��·�oS� J�)f�\�D(#�B���Wo󶝹,��
K���u�!cϓ�� ��L��4��y_���� ;�0�-H�c#�ԃ�ˍ��~��D'I��t���Yu�'�.x �{�y��AW�C�L���V�3���	�^�ҙ^����I��a���� x)"4NqR�q{���!n�I*\ᥩB�=4�.bk{��t�O 8��ɥe�H�(A�� `��i��o��[�֒F����-%��;�����ā��B;D����p!]s�y���̀�G��9f��UFg�u�Y��37_�����.¿6ep=��x���Q����d�����x�SA.9���W!�n�L��.�	�I�}l�����CZ�UD��J��ZQ[1�Z4��8��pi9�|�#�=�(����"!ri>��9�S���v��ț)��ʓ#<���B�|�uj�0ݷ���%�>�@�:���d{=��`l.�CF�^y}�XTOؘc�6m<_��~��J��d	�l_2����Aytё'!��Un��E��쾥�%Nb�ȁ+֟�<R���)�+_gn���%�W��k����侼R�y��+�x�#+�������.��F,{���|軿�N�\X�Y���i�һ��Z!��p�1< ��/���0je�~������i���'�_���u�TT>Y�D�ꍉtv���Ԃ�/<aG��*�!�ք�DH��L�Oy��`d�
+�����Wɩh!o���(p�=7K�
�}�*���U������rT��tS� ,�sA����_�k�C��3ZI���Ҝ�J��]��z�;�.<�_>��AesdU�����2 ��H!�\��5�1�B�'o��z'nr����+��@#�m�[����fA��/�*�a8���dOE�K7��0,��z���^�i���w�f#��A]�Ja�\��
P�IȮ|A�[�pIl�au}��v {�Ay�"Cn�=�uT_�����
����JkK\+*I��B�[Ds�W9�~�C���$nA1�5�oG����=�
��vα��W�;�>�bZ�v���7yx��3E�oA?D�z~����vt�����L=?�	�<�(�ΐ�'�ڑ��!@3���q��}r��G��@��ĥ�0����V*��sUIB5aShe�piʔi�G�<��[/p�G��z#G]�G6���j����XON��ӏ��d��R4�Ro1��:u��q���5K��Re*f�W�]��Y�ʐ#d��ft�g����9҅�B����'1y�h7m�'Ac�����_�4�6�k|�k�O������ ���=
֕��E"��)��h`���å�-��G����0�-���a��T-0�������#�QL16�\((����# ��C��2`���� ��\�C/6Z6mި�E6;�]��o����ۛ,n�$���{Q#;�K�H�Kᡣ�j#�J��$�"�
��{Ȍ��̡�;n�H����Ř���e(�7��}��p(���X�)���jV�N����°X56�u�HB�Z1�Y��͇f̚�.�����mג���i�fc[��?�c�!�>F@��:j���s�@�)����̌6;V�7GG�J܉T�r�����%B7�Y@Gjԏϟ�%�|�|G�G;���1�g6$,��l�Gdd���DB*G2�5X�U�	rѲ7��J4�vy��M��#��3�|�RK/$Mf��S\q�LRPA��UkU����`�;��2"X��Ƭ�Y�-��g��Oi��8�\%�������q뻂�b��X�y��Fռ�PT�e.\:�v\+v<���]J'��C�I�^a�dO-���O���bt�<�$�ǀBg�t�I�����KC>Oh@�������P��爎눎瘎�J���X,���fWԲ�2gv�v���ѽQ�������3��`��
_eh/=�%���rՍ�ԗ�	s���:����Owع����(ȷ�e�T�t"�7�|�������dqx� ��xC��s:�hA��OiI����5&UV��አjo1ݮ��^	�m�S)�q���Y�*kk����A>�n�^\b��o�o �$�5���M�#��o�Z�i�J��**J� L��Uǯa�PH3�vSM��n(��I����F���]����$D�*:9�o�{O'���'�te:�<h�Z!Na�8�������(�q|�e��+?E2�0��;����8D�&ozm'Q���l�$�:$�X��>S 3؈4�{m=ۤ��a����c�b x�>"�C\��Sz��}����ꤑD3_�	�9�Ă@Br����`y��vI;*�A�w�/��6���w�NiYŀB��=��C�kQz��Qb�Y<?4�R�=@eql�՟�G#�W�f��`�-900+��T�%�D	�������I�=�LŜ)r�T0q3@g���DD���
�~����*Z����S%����Y�UF@�q++������p�fK��}�/�,Z�ւ�Ǉ
���<g��L��p�M_н�Q8���C �+ֳ�3�S�$r�@�%���Lਹ|���h
������i�a]�j	�JȐ%%�;���N2m��!���dXhhp��C��M��ޙH�#�w��l�{�k�cJ�3-�1�y�,�qa�zL�T/��b�G��ܢ|�M;gob`��SE�S�!_�m)\�1����l�m�lB>��u��h����\B�zAT�cZ�W����e�::��'cCC�����]J�{u%������'�01'�"k�����\!ބ
���׆jG�B"�9�C�@(&1%k~l���C|��*��� .�R���k}�PڔD�J�5�M�k��E�eY�����U;"�OD����1�6�Ep���Y�G�8��Q�ZB�`��A�m��̯x� �I1�1��9�����U���jD���7�ޙ0�S�Y��i�yL\;;��V�:!�Օ(h�aE'fs��*;��Cz(�Y�KBV���"*��:^�ڲ	Xጂ���z^R��Ĝгg�߉��3YW�F-����}!�u��B���I����e�||�y\A�B�.=ՉS�� ��-���zH_���8���wևNIGhꚚ�-b"���Q���f7Zl�=لYnY.�V���'[ �Ic�>���s>q��"��w�믨׈�'�6ۗMXdQ�%�f�9(>��}�ɘ+H��z\�O�$��x���6���~c�&!c�8H�0�1�I�ҕ�Uzp7�l�]8[���]�����60^;���]FQL�Q����d��A`�w�8�I!5�:
�^�[v�XV�[�#��!�4�T�ɲ�"۳2I�!�h
�X~X�7�?h���NǮ|���o y#��4�0��t߮*�6~��
{f�S�����$���������׼9�L&�A3U`�Ȑ�'�$�}�)٩��H(�tL�ژG���@,��'Թ+�*&5�Ӫ��ט�y;,d�.�Z+VB�0����NR}�&E�,	�O�6z���^[���ca*n�h~7gk�߰�O���/���cd�-�
���S-��V�_B��#U���ǀ�=�kO����|�WM�
���qV�n�5Ò|�ȼ_g��M��uֲS$����`���:���)+��3�P�Q�`��]�o�^uӈ��ӸJ��9G��|	�IH���jH#����ru�W��I^�H²�T��������\)r������^!KT�# �y��gtT�L�l(�����Pn���5Y s������vp���~
��ߍD� �e�6�j3 ��!H1��K:����B��o��Hi1�8�"x�fRЂ���j�l!}H��c����F��.��ԟCr<��!��9PQ?!��r��q�#"N��-������_G #���NU�dK�2��7����Z�:BTh�Qj����^�. &���ջ�<4:����<���uZ!�_'�^��^�k�/3�)*ۻ�E ���lb�ζ*"岗����f�檱܃x ���Ude ��t��ğ[~?�ڹt�:U�o��ؤE���9;\F����UQf
x��*L�?�^�w��6��.�Fa*�W-��T�V�.Qj����^���D{��j��ڸc}� 1Kj͠߸�D˃^�{U�0>��B�Ǌu��������=Y������ɶp�����;C�!�&Ls��^��L������6����^�2����4\^�l�`�ꎊeB
�_���I9�#�;+�c4����F�XH'����k�R`��g��;�zt���n���tF{ׅB@0�^�]�.��#�4������ƴ�� lM����b9%!&J ��\#�j�����do �i?��~P��/<{�.Qh$�CH&b@�����!ϼ}EYd�qK����}x#e\���d���!5 �q̫��V١(d#@9Ś1���)�fqU�	���_�r,�C�]R�T��Be\���o/��Y�Z�dk��F�4!e�o�ו��NB[��Ql�g�U��7���f�W�`)TkfI��(JW2�1����1��'䰢k�Ȣb�n ����%�g�����Z+��m)��&�;�E-��-��Z�I��mD�0KQ�.r%.R�v������C�-g�A�k|�@�r��8k\�ՠ�����I�au{i�]��]�]��z�M�@�?kF`����w b>6Z�(U��c����@ �d�R�H��a�.������:�s
ѥh�Ȱ"I"��p�4Ȯ�F���	(���摨u@B����wJR�p"`þ�@�T��PxBE�����|�=P��N�@wx����³Q�_�k�TI���_&�/~Y3M����_�ƯE@�U(�녉
m��D��D��m����,6�w% Lwt�_ɤr4Y����s/��nN*s<�N��2 ���P����"j�<�t�	��8��d����b��!6�7N�@��{�P�Mc#VHT��Nk[^�y!��2jw�P���o@�j�&9\���J����&���)�x�~g(�F�a�{����RwUHL/��Ф��������G��G��PI	�$låJs/^�'�I{���B3�����4����r�Qܳ!�V)�h)�B�-;�-�#>���l��R�@aZ�B�ut���T�x��p�#r7l��.͐PG\�G���Y�<C���~~�ϱDV�^�kזР�d�'/{N�hs�Iݧ��2���v��RMt�-2af��#�s���F	�S���25�-M@���\��7N3��>���䄯ͼ�b%t���3q7��/6pg�I-�徘!+�.��j2ey��G�U����%�G �5U��"
R(r'Q/9�?@�(IVI&D���3Z��iⓎ�zc�e�A!ޤ�W�o*������A�ʙ{\�T�?�[��o��I"���{4���odO��i�Q��.�<)�f�x����-y+$J6���Q�)��LN�I�QK��Y�D�=D�fkR�T~jv T��idL�1�TYr�vJ5��D q2�����t����I�R�Tj+�;oq3�҇CA�4L�#E�]��J�x8�y���l%��سR� y'}�H����)+�������+��:7W�$�">���H���N_��|s���W��Cb���Ϣ(�/)�=��]�@PvF�"�B;K��ӻny��D�����^FQ�2�Ϣk�����'ozזkR����Τz�{濫��h���<�}�8�[�L���3���m~l9�;)N���YbZ�d��8;���^��/�m��h�/�yu��J�k:h��&�x`�!��[�E�US<�.0�o��@@���tx�=�]kXC��i�m'�T#�z/9؉6��#	�*Q5g7%���|b�?"iE#�%�e��v�
B�d���m;��qv�rY�䛇�����DL)���C�[�E�}Q�Xt7HJ#%-()�tK��0��� ��H��-�Cw3t0�>��{�?���>��Zk�s�KX�$��HTg���y����0������9BJ�;�s��3X�w?�T8�d��\(��-a�D�LO�o!�O���/�C���M�1�8{/�L�;���&D����Ǫ��W:���UBBÍi
�)�H���dT@��Ǉk����[�=��ZX�Cm:�JS�(_�G���u���i�N��f������w˒��)���cX�v�a��YP���	��'��?oR��Z~�p�	o���4��i݈ꢞ���<�����] ���գ{��+�鞸qO�i��^,�c2{'|B�rL�����ǲ��d���
Y�G�����$�� �b�S
p���畉p�n�[�O˭�Xq�[_@c�J��f@��T��_�y\��Xe����v|g{�%��Q���Q���-+��e:sβ��R�ܷo��h�{��1��E�����t@4c�e֊ ���P�r_Y�Y��swm����U}ٲ\o��6O8�\E�E\��M�����T�e��u�}�ߠj���b�f�#��_�;8콄6�䜙�ˬ�>}����G�h�u��pzU�<��M�y���2v��P�&#����s��0Q�9a4#�D:�Kj���������W���N�>���!I�/�S�ѕx�]6jű)	�)~8����(s[��.�Qu����5 ��C��>�_�r�x�&�%U?�E"�4��#�X�pf[��h�~��i<�Q�8�X��L���a;�P�ebz��l^ͧ�>�����Q��~��B-5>7s�*�K����񰤻V)~���S�c�:ߧ�q=ky�5h�W)��d�½��4����������B� �r�sӹ@��r�i9	���H�����W��$ؙe^ę���E�Źs��-�3�2�	�6{��_��u����G�s�s��߅rH8��c;�5)r�+r�� +�i�����/0�y�9ʹ"����5���5�\.\���@�g�1�^l2ʣ�;{�Qf���>a�	2�@������hW�����H�Fnވ �|q*:�}/����͜��d�h�\h�;G(B��u�f�)��,����/k���`����	?��o�}�:����6�9܆ ����eM�=�|��O!���Y�M��~~qQ�[P�{��9��,|�k�V�x�v�AT��0H\�L>�`)��Aѫ��;	Uup�^څ��eoбa} x���9����B9ϓ�Z����
?�0A� 1�M�\U����7Ek��9lnm=uΞݮ4�t@���ɾ?R�`�%��r�s֏D��5(o�>��� |ڗ�Xq�>���yI�D ��O; Ҫ*K��Gg�� ����G�"7%b��`�1�-�'O���d
�u���{0ZNZwO3j�[=Uy�췥O�� ���e:)h�aST_<�	�k��+�bK6�:�3��X� ���7�(��!�Z�d���i
N��N�M��퍽�ّ�є����]�%G���=a��z�i�Љg�J�kQtBg�G��z�7�%b:[+<L��b�3uu��ޑ.�Ћ{@_�Ϊ���dw:�V5R�/�duq0�lC��&�!(�I��X
W��:<���&��F��$�W�#���p�T��)R<B�j�ծ�u�k-�n���[�S�Tě���f�6���������X��遨�_`�¥�ө����0��Ƕ�%C��,�V��=�j�۴�TCu{�����]�.��f������vZ�M�IvAԈ�^�A��=�J�;!���ug��w�cO5����殍��Ϟ���Jn�*N�)��쮢ff�_�S��*�W��.�Wʘ�Y��d�L!nS�ƪO�FKo,C��aLQl�a�Of�b�`��$��zZ+>tB~�l- >	a��ޗo6��0\�`cDz�]���B��]�F0&JRc�j�Ԣ��h1���z���U��#�w,��}�Y��d�o￐T�5<dy�X��-�&�hh$����h�y
��f3LU�����W�U~�ȔiDܮ�h�l�9��d4L�:�g=�z4똠����f�[y�0��1�T��Uh�*7o�]x�`�'D�ޘY*f����S=ܻ�T&�;������J��C 
yO):�Ϯco�`q��)�"1��$
^��uҡ�B�^��u���qyYĶ����BѼ-���&��;u��$�h�]T�s�d���b�Q���D�����3ۈW����	��uz���k
��z�lū��d�;���0p�/����,DہyB"��)���<G��fc㜡7�a�Ki���#s�O���(�� ��Х'�p{]�ȭ�y+Z��O�����^�l���Z���|'�p�[V&��0�鳶.*bleBx*�����'���x�_|�IG���ӑ	Vf���p�t�+��3�`�`O�.���@:�����ϫ�Y���&��gqz�C=L��5�#�m�b�K�&,�^y��f}� 񈘏� D���4)Hx�otS�|=��v7nӼ��5R$�p�{�t�F���@O�뼆�(Q�mbv�'�	Jl����	%�]2d��bƟ�|�	H3��^;(s+6�wطX������$զ��|e�>�n�XS������5���
��s�$�x���MCG]���nN 	���#�ڲ�#��$�����S���N�4Kp���tr�h8�Rh��2�)�^��wSk3(�Q�y���m�����-��Lr[4���m����ş��k��܁������Y � B���ݡ�N/�oJ�6Z.Ƞ��ƽ$f.�?��j<+�kT��6z�҈:KnKޠ��)
�6y�m����W���ʹ��=}�C2��Wר(Z��ՑN�M��dO�F,�`�L#�����G������/�����tK��E�	�vF:/ȏ9�����J*i;m��6�s����ڗ����)�=x�����E��f�PEٖ�����"���۫M$L�~�Y��{�g�~@9�@�������$d�#���;�Ki�̒:Q1J�x.K�ܩ��f�n���SO�&���TB�E��t���R�5%�H^�1�6Wd�U�j� )c,�s��|&N��<=�,�1���K����=�}�z�)?��Y�.9�%�M��f4 �E��j����x� =A�_�3&!/3V�+�I�y=ڢ�� �ɆJ�U�{.Wd57�5��3�����U�8���e6Y�#����gWBc���|=���������[�c����yAC\:�l��|���ny�.1��� ��u���� �^E=��ٹ��d%�1*:�}鿫���T��Z���b���kҥZ K�7�N�V��b����at���W��K�篧��˚��J�y��
���+�.�����"^V�ۧ�5r�K��F� ac�:��O9�M�F)l��l�7��~�³�����?m"���^P+�.�{N�qe��bF>�kI �V��/��?)�R�^>�@�7bgRA��8x(����B���Y���P����cYʊTp��Zn�%���+
&��t�1ōh4���!�h��a�j�Hŵd̐M�G�y����V1���!���7OZ�vv��ꛏ�D���Ku���W�;DV��uFM:��~�P� 8!)^tjF8����:6.C��g��0��&�R�T�Dw��#~�<B�_-�g^Q��]�3�RK�V��C���F���$����I�Zْ_�4��E�;��z������Tn�����@��>AK#�s��,i�����X��$�Epػ*�s��(�m�) �!ϣF.~?1�]Rh�_�U!�Ev;3���|�� Cݯb��_���o��)���흀Yi�;@�{��2�z�>y�Ө���׌�)K���f>Hb�3J� ��B�V5�����!�_Uþ�S(g��˒^�&��{����F�^�U���z�AC�1��Vm�<;M
��.6'����>�@Eބ�;{�z�$P�RnCͮ��+{6�O��WnR����5���tכr����}z�5qV�+X�2��ٷ
~5�$h��%���m�9H�Q�[����򣃁 "�uGЙΓЊe^�^-(���!��j䕋m�W#�}-������5z��"$�X߳Iګ~Z[�n
hW>7��-��_��߮��Ү��V���w9�0t�ӟ��Tt(����L��;�A�lH�KfV= ��[
��2��K��-�P��b��U��}ӷ�.�����D�\�y<�tq�Q􏃅hyц%��o�ރ�n73�6Yi��ʴ6��ܣ��R�So ��b��7��ĊTM#z�:f�	��ԝ��ˀB^&Վ];���y+$eTv=����yֹ^�7����[��KL"'Ϊ�������O��/RW
L�hﳬ�Z�j�D��h%JHm�娼��/�Vt��ndV:-��Xi.�i8���5a2��`���ƧY�)�����bq�v٪���TZ[�k'q9B	��͘�bY��B&l1U��Cc����PM	A�-����©�&�'�˪�۬PW�x]��8$�8È�e�*0�Z�����oo����;%�3�K	bk2c�o��r?�	�7x���T�S�	w���CP� ܁{���⵭G ��Q�Y�8}���ΰ����EGIź��bd̗l�u{����k����Kl�!)mR;
0�r�I%�>����N'�1�u���Ԝ2�+Q��s�<�ed��GY� ��a��8���#)��$WD��`ư����L����I=�j�.��3�B���(=?�B�+�ܹ�a}V��MrSn����ϫӆ�}�+C�_d[}$;Ӏ�:�r��`�#�(�[?E�o8����3K:�T�;$��}���g���Dg�Z��r���.�#<by�����0���8�C�OQ�u'��@���W;$���43�t��]�i�N�g����5��� �oz�d���^�eV��lL���Wo���HCO������~[In��Z�G��#�ETt>�
�;�k���ּ���(~X����|�\�H�w�E����8���-���v�ؓaVrFx�v�b'p�*�0��㗧ybYV��|�����H�J�i�L]�v��.��#�U����%�b�� ���E��.���R��(��x�)�{�����3�����m���EQ��z�P4�^̓r�\!,1վ�

�`�X���'����B��z���Yt�-�Et���Η���F�y�l��>���I/��r�Z�Ia�yf�H�^�u��d �|JE��1h6�
"G���?��l����z�I�	�u��z����t��<*�	�t�9��q^�O�Xe����W8�90��n~���zeA�0I|��eg���3��[�����Bi�&�W����cU\��	�#��9n�"�C��q�[d�7Y��K-�hB�-�:����y-T�V�s��Z�c��Gv���g�A�|���%vЉ��`B'���o?9�c!O�Zg�^SsNb�<�rTk�ٯj�ܴ%���ޤ��/k�
�P���M/��ק��+����G$��40����O�{ʼ:C˴����(���2��9��[�t'�{��\F�ot��H�$̝�Oo�긏
6�g��=u)����xJ���(iVS�
Q#��S��g�i�]��8�b�M���"���:���l��������ي��|׫�i�jTF�]2�O~ױ�����"h�o�	�v�n���R�"�?�8~�������>���~�ޗ뢗�AO%��y��\���R����nx6�vl�� �0IR��|"3|3�.՛�CR�\�o�Ʌ���v�Sx�V*�N����'C(�:�{0��#�%[�#s1:�ヂ�6�cL�h9Z��?8��ޘ���ֵ��-�?|�d�mpR�p�_)��5�37���ƥ��m^+�ܹ�s9��7�?�'^��ɂ�p�����D��>y5�)	.Iwk�kKn�K�KlsBI f]dG�9�-���HﲳԎ���]]�O9�*W{y4�:61~2�L�ī�3���ߤ������J	���c4�Y���&E��Y�*m xH)h,�;��?�K!���x.Zk�5�K��T���\&�J!Ixc,�,��;�l�C�&c��A�b$`���|��<����&9�nk6ۈ�&��g唙{L�LAa��5Ɠ�U�D� ���l�b���D��"�K����o�i�҅zN~��-3�חq�[�H�I�&�v!���6T�I��]d�O}	޳>�P�FD!�����A|��So߸��ȟ��Zŵ�\l9(�M�g�� ���d�7��)�i�[�0'm�pt?�*�� �`"��QZ��@	�Ʉߥ��(%D)F��W����oA�+�q�_7G�xd�;mVīNgԚ���e��:�܅��:�֪�o��S�;dN�}�G�|(���F�n�!�q���ef���is�񜵧��:����S��k�⼭S~�6p��h����W��i_��LUT��w�MS�Ȁ�������R�.��
�BF���]5ԫ��U?g�����K ���<�Z{�]d��}�V�kσ��T@��2�����?��B���>�|~��r���?��ә��s.9Ó/=/�/�
�a���Ήp�X��:�Յ�jll��.�<�ܳ�!�.�"l���-[s�j�n���:��s�������O�8��3Սႇ�k�6ǰt��X���&J�b,�[�W���SP������e���9���OÊz���t?d�U��T/Va]�s9�B\e�	��bI�UQ&�Wm3(� M�ۉ�������Έ�����*�z�2\hf=��2!*��}��_�x�ڠ�;:W��"��i�l��e?��KG������e2�Xg�6�ݮ?��}�p��E.��1����%���[��i� ظ)Z����V!�tc�e�<�7,*!�s19p!���q��α�p��p������|��K\iǳ��=��h!I�_���c"�
���h��H�z�޻��YR�����l�}�[�"��t���	�%Wq��3Rf�����X�zq�9�5��	����/Ua"�}ڵ3_ׄg��:39'��_n�F߾�NS�)����ij�gU�{Dr����M�l~9��?�����&Z�|S������*���W���}����YEH���<}���~# w�	A�%);Fm٩Ȳ�i�����{��3�+���ܭf�&����-�X���{���+B���~��f�PlWC �#i�O�`���?���p��e����j�+��M!�n�6+��2˖����9������\K�)d�e|�!FH!���u��"�ip�e���x@���g��ڧ�I�q!y7e�ޥQ�WE�+C�-��v�6��T�8��zb�hMD�Նy��|�(� ���0i$<I0/�r��$J���8��ٌ>�R�[M2�i��y����~H�\�F�PQ����������>�$�X�,tM0�	��n��G��0��[�HI����r��J��"�̿H;ȡ���ķe¤�*M/�_03��%J�>�o""��vȜW�V���AP���� ə�űߩ$x�B�6 ����WД.nۡ&0')K�ӕ�
�$Z��K�t����J?�A���w��&G������<� ���Y
� �ÿj��@� �����;��G�pďqc:�̉ƅ�l��V��iv+������Ռ��������
\�Sau�3�.�!~d������S�B�]'�G���,��4�sH�ď�`�s�ml��SP!�i��'yynU���]`�[��������)��D���r���W��yl3!K��!��Fq�r����b���ݝ�T�m<��>�GuҨ�g}��V�'�H��q٤}�3]�\�ĲyEݛז�!I�s�	O؍q�%�h���Zr�V�=/�Ns��1�.l;=�2��d����㌷m��L[�?��ꑬn�Kw�IP	�RBü�md9����x{��&�w�-��)�؆V&�"�#{�j�%ܤ��l>��$�tz<Sm��H �x�~\"�Ka{�����5���ܯ��%My9��ʹ�=�����m鑋�4[��WG����������<�3�d�Gnk[)R(���k�s���[�~͒��8���-�a�
 %��j �5?:���$!l"�z�myv�˞�>y�']�xT�v��lţ6��L31%�bC*F��Y�=M�.VS���xN�*���%�%��}B��2� ���M�7[mW��T�B� CQ�㖅�&�hrW��D�.z~U�{�e���tF3u��'��xaTM3%���+����Sr�b­�^"���y�k�`%�z]�H�a�]���Wm��8&H�Wg�O$XxM�7��p\(i��v�ےfS�s��|\qHN����gc���v���Y�9����<��1k�x/1��d��a�un���3��y>�_�j��"��h�0Gl���8�U���.w�y��NA�Ŗ� �����h?k��z=��̘H��������Mr�4�v �޻�v��{��T��G6[���������8nv�=�
�c�V$}��P��������ӛ�R���W�Ѧ_"�lD���a_�ۥ9�M��c��)2M��q�VH��� `3�� ���*c�&�' de��+3�-��Ρq��� I�1.6�M�r�gd�N�4�>���5{��8'8�t�۟n��%ya�O9��eT��I�42�P�\ke���~������8�nC�Q{-~"R� )�C`��(��2,	圯��y��*����\��F�J2���r��}�'�]q�l�ֵ~�����K�X��t��e�'D.p 0�#��du�8Imn���	(r��'J��I���g,H2W@E/5��qȂP.��>"�о���*{�pJ��4^C��K�0u=����IHa@������\俰�x8��;i6�|%x�5V̭���h��F.��[o��M��%�mc	5[�8���6hH	���2�$��X7f�Tr5 ��i�F��9�C`���n�����vb�c���y�re5���~���7:=�s�FH��p3ǔ=־��"Hm� �ԃ<��=��lX�Y�pL����o�`�C�=or�M�blU{=Iu�<ֻd"(��>i��]���H����.1,Dї��9�B�Ӏ=nQ��A/�ظ���f���R_�a}���T_��{B����1�G���R|K\�d�f���	���t(c#�� b��*G��]}�'U�~>Kҩ%���w�r�s8��q
a�i����CҮuQ�*/�����k|m��+���^O/k����xy�x�w��`��=Z�)�����Χ�-w����_��k�8��'d���ujiW��}���C���������í*�K�+DQ�������3���R5�<�rF���V��_�f����倲Y�������D�o�<�̳`��GrC��+���2+U�Ƿ�[?��x��m>�e�+�|�P��c{F�3��f"���8���tji��&�޻F����}B~�+_X��T��f�i�/�4��?�D,d��>���n:7i
ӫ���m��ִK���q��3���Z�.2�hu��y����`(c��W���ݶ�ߜ����|��>��5�ඁ _*B'= 5s��I-is�nF�Bn��	I���1GG��Wl�ƁI�7�E��0c�{wf��u�u��	�C+<�{��v�����k����9e���-&s���~(�FʹI����$�_K��@���=�5����Ls/���Z�)쫦�U�}a�
^��-��2�Lٳ��@����wz�ę�[�~�h�.hA�Vt��4�7�P�������Ϋ5!�3�����q�@44��)�� ��<�oC��i�I/w���Q���c[L�	����M{W��^i�9�rLW�Y�|�T�ۄ|�� |��us�+J/bh%�QN��Ba�/�aD��Q.81M�S��Y��"V���/�X�M/�����
����KF�hy������ ���hN��W�\�H���`��1�Na�����������n�@6�8��5�7؁~XF(�i��d��{̏I�M�����Te����{���jG-��+ �F#{�5��Ch��w��OE����o]��/���L.5AdX�9�����g�Sg��Nٞ�nce���F�A��4��t����Wyw���N�;����x0�u#�:�N�ڲ%���Ѯ��97�h�)�Pr
�K8�TUТ�+RCsV�/��LW��Ɠ�4�X�\��ڻu�l%]�5�®ʹ��~n���ƼΦ�R:�h�DiR�gÚ��_ƕm�t�^胊�Rs���:�H��g��L�+,���c%t.k�)c;�	� �͒�[��������+A�E�9���h���`pV�D�4}�Յ2�ALX\* >̌IB�M�3��p�Ŧ]T���5q5
�vӊ�T���Fv>����v�B,��M�ҙ�K���鶽ܘ|8�4�hG�M.�u�k2G�b�v�c�:�]���hȯv��9��G���P�^ԍ�cE~&ʓ�mS4�OT��6�2��Av���������)����!(O2-\�Nb:k��y��H�����y*x�yG4|oy��7�sݟt�����TƐ�z�B�y���$(���t���OR����]��GH��~f���;�`ΕVM���!�|H�\�Wn��Z�'�^Һ%�X>�.p�����Z�zm��eN���#q����.��~l��Ua]�P�r���	|��SZ;rW֗I;��}d���!a��R�kh-�՛�1/	�B��]�7%�ll��b��dI�@V��@vKESO+��Tm�}�k)�Ȱ���qͣ�q茌�VS�B<�\���R/���qD��ˉ�Ӻ�ڽ��E;��z����Q3���	 ��`�-��/��T"YZ��G![���L4�z��ѿ��a�7�-5�X��%: �t��l"H|��p�_Tp�t�'w.��l�Ye���C0�3:������E��;�Y��z����_�XN���u>��5v��C��_�k�:by��g����+��L[>�zn,l����$z���t�N�+}�0L�0�+���F�t����u�!\���tm�B)n�Jebe�߄�.�|*x�N��n���z"rHUbNT�i�;U5�����xG�-�w����m���I�����7��e����O�9�M�	�F�<6�ŗ\�Ҧ�)�!Iب�Ô���C�|�]�
�;��E���;��D+��95d������n���318�ihO��͒�pR:?�5-�k��6*禝$�Vnв�$��_tn�����q�*��p���r$Y��R�"��ˊ�U3����5�Q
_��X���9�+���	p\�p��$~��E	Wnyԛ��l�yS$~�~"/�aȰ��?��Dʶ�8]���FB��=6V ��� ���k��;����g��3i�4�0Q�>^?R�s��l����p��bf�vپ�p���u$	���:v�q�W����5)p�|����m;�2����>�_�4ꍦ�n8�]��S_���v��Q�U6G1R*y��c޸�	p>j�Q摒T\��8PGE�a��xϬ/R�c��	C��U4K1*bs�ǡH	��.��Ѻ�G�Ϥ/Hq�]��"��X�]����I��Ӓ���0�7�b6~��SBI7Q&>s��ӕxs$L�_��������c���,��Z�7$��ڥ��twM"#�b��;�q0D֡�dd������s��4�'��R�2/i�co����o����G�!�^��^Tjl15��`�����u��b�	ɯ������g��	+���1��>���/3�w_
��E��2%P���_�q���pw��������up���,�g��� ���CJ�.�:�j�<��ʀ�k�m�ӁԎ�)�k�q���h��m���%�:_,��p��'y��?N�t��)Mpm�e�[̇�_��>@�*76�b��&��l�I�m���5���u�8?i�����	/�%1���9Tz��`0��|
�Hk�2g6�떦��c�x������������ϞM̏dCx2v.[2�ZL3׶Cp.��Fht����^aY�>�A����w� �s���V��͙��s��R�asc
'�nL5�N�c��8��ςL����#��FS�^}����P��U�;=�;9=����2��B/��/�0b$�԰˒n��q�|$~/�N��qY9�%io1``ȍVR��X��y�Ȥ<�䖇�I��ŵ�n�
�c�i�:T3y��į�r�,Z�,�����LJ[��R;��l����M�E�ɡ��-ٮ�~�},���i�g�4�?f���|p?�whW�k�'��wŲ���><v�s�u�+������������CfЦp��{np��#��IaR�O+&����%�D��6ϖ�
��w[գ�+���N"{�lP�ӱS�g�Y�D�|���P2yӔ�]#�n��+s3�b���+��*��
�X��m?�O[�<�o�6��j:�!�&��k��z!��Q'�D�_�2�>))+Af��B]t>+kd����"J�3��3��$�z�A�+�lc��o}�X���e���ZV�x� iOqhT-A�$�ֿ�s3�����9#Zh�>���x/�8���p��3n�"tB�Fn�p� h��ئ�6ȼe�M�3E�r���/�w�k���y�/ Q�sڟؖG�9���/���4����&��Y�j6�fa\�؏N+��߿��JOv@��B�q~���y���쁉� ƀ㦒���ꐒ��N�f��>T�ȀmhV�s,�<�� �6�Mew��%��Y�����Ʒx�|��k���7�ژ����R����g]�q�����|~�P�]����$�^�E��{k��o*���A�R��ɗ�W�R����#��Do7��<�8"�$��8���}���\��>��L��rlߑ���s2<N�n��kV��(�j�
d�x;)bR�%1�>������&���!T)�f<�P�j�7tq�xK�ejp�i��2N�l{:�	����R����vH�a���i�Rqpk_���X`�-nfi�c�a,�	��<��.�쳽��=oK#�?_��4�T�����@o���zS8�qǭ�f����4%�KϺ��O,���a�� n�Fu���"鉊�:X��V��_L>p4m�˜é�L_i��!�"�[��ɛ}i���r5�IC�NM��{)MS�����e].F�r���hh6��$�f����f��z�3uE��j�YQ~J���+�*w$�������������uvq��0���<��Od;N�-x��x�/��	��;�ܙq=�6Dy�����mv �����(��T{jO�4�/W��]���K;��Un�l}#���	��S����-����V��MdC����;�Y��o�
�Uun�(��:����c�?3���s�5�[ʋ\Ba�'���i(�C޷5�̂i���?W��L�OBᗙ��t��,�ݟ@K>�޿���)����^c��%�VvoVG���,��]b�����x ���|���8�kC����Q"�I���=oɰh��{�dj�֮�(�r�h3�&����vb���U�㛎S��#��7@�ѩi"�5"������9Ξ>���(�5mo-��<���6#*u��2ތS��z�%]��q�}�	���~5����+^<h=}����|�O2SP3*�!S��d��r�RR=k�V�c�Q��hk`��f���fq@��et���p��F�6�V�n����X��K�v��0��e���e�A��Gq#WB�Io1�cv}��:�k�6��n�Ȼ-��E��\��PEŕH]�oL��3���G)��m�V�uW���Co�k���b� ���TW��ɿ���ıK�.p�4n}'��@��������T��wu�8�7��f|F�qn�r\z{:I�h<l�����|��]����@N-�I�f�>�mbu�kq"�Z�A�"U|���I[��&
6f�����?2`��PB�D�tx_�YS�`�%����D�G�|���3��2��򋕹�xW�(N����m��\2�=.��>����3���Lq�s�)m
�j��X�՝˚��Z��hA#�x3�\��I)�19��3��.�J�af���3��	ق�aMF��4��a��T��-�aY'r�c$�s�£߸Atߞ7~��'_����W_$&l<��v����c��f�ӊ�t</��KRF��m��O��<䕊B%�2$Pj��o:uڧD������,�1�S�+�{}�	��
��R���r<`�J����~� z{������*�969�iU������Y�d�}�?��I4�� �U,H�k�i�ژv_T�^��2FjI�����>�@�]3j]�}�z���"�Wq�V>�4��E>f�m�
�czV�"쀳�'�u[�}ékgG=�O�Z�³��&g?>��:�yJl4�m�pP�6u�B�ym�My0��}�0�ۍ�'�a�ϓ�W�mpIɣ=��R�b��fmt3}���w܈�Y�2�	;fYP�KYü�!�OY�I�b.�����g��jY��l���ni<q]��ƛ�����Zؗ�u�z*���`��c'(`�ʷ�o�#�aY�	�V�I���������%&��E��g�f�"�w�p'����5[�	�/�;�R�I�3��2f�7@)��j�>;3
�xލ4�����<_��#��XA��kS�C�d���R�e�Xl�H~&��-����QA��e׻QP�>0�xϡߺ�x]�a�.��P|��H_R�ae�z��pe�S��6K���x��la8���6�&��X���%WL*T���%_�+����}��ղ,��A�!f"ʾ
E�����T86��>���N�*�0�:kh�D�]�(D
��i�Ƚ_�n?}��r�/� ]�W�f=p��鉇��{�\��
G�/b��}wgE��+1JӘ����|�2J�L3n��#������a��j��sY�
pd��������0𮂾ˌ8�e5=�j��7�>�,D� gї{���N����ў�A�z>`�rdt����(�@���ƞ�D�K�ޥҶ��G���<���$s����5.���v�ݝ�R>9Ȫ���g��g��c���)�6$�E���|�h��z���!$����<z���l����4�ı��#|�����S�m���Q�/�4�_�ʜ���l��\Ĉ�k�}j<iik���R�1<#��ux]o��=�͆Ȼ�B�:%9h���������-��By�oR��U�-����<�ł��P�-�ȗ��j��0�����ȍrׇ�ذ9-�K�}M���R���'Q�3����/��򂣓��8Mz��]7QF�s�V�]�>S��z� �'���^��4 ?I��/��?U�,/��L���n�`�����|�REy-_��9^��Fuݓ��E�*A��k�V6ԕ�Zib�b0���ҭ�4|�����+��u��W4ft�L1�]Gv�}�]p�[�R	��� ��v��6˨=���ZH��>5�&��������B�v�d�Ƀ1|���elmB!��\$t�eM���������^�G�Ԑ���
��:�.�zG*�Z��dm��e����^��p��e���F���c�s�קM�=��|���>;" ��?�15P� x�./>$�����8��
�6���s*X��)��u[�zGc����B?U��C�?7d,O�k�{��N��;R�]{7EՈ�2Ծ��b��P�y����ȧ��ɏ��g1�ы�e�j+|o�i�2�#�I�r_6�#�Wh����*>OuF�%#��k09����P.��`)ީ� ��3���f�(���*ڮ���!���+�&	y|���3yD�!p1��݉��M�P)���U�3jwP^���K��-�0@d�UvY�q� �!�&F�h�\��e��	A}�&D���?d��#�f�}J�㖬��Q��A��Z2B�Xd���=��X�I���Qrw�]�+��<`s6�?�l#��:r�O\�o���_����T��F��sg���w;k9��!���)�~J"�Đ�CU7{�A@���nv�&ew�L�+R�7��Ih����F$�� ���w�y���@ Lj�dk61Q����a��B�}�L�|ki�.1��M1
��+x ҅n� �H1���@�n6��F;����b���<��m���s�hBL������
�o�$ �y�2G���������y
Q!#,�n)�U
t�_�k'd��}��pF��O��I�3��t�?��>� Z�H�7����)�/]�}B�&���H�?��
�@x�P�;t�i�u=��ox�՝*����?br����&&�{vOJ�UF�x.�v��Y�c����
�G�##��! :�Ț�Dп%y�G|�=��{4����s�Z�AN���N#
i �����%c���O��]�S,�"�X���5�Z.�y��ڥ_J"��U$拏U;���L���= "���J4�GE�M���<�S//˅�~tm��TM��ٍ�/^x��*}�5�Cs�r��)���o�8��U:�p[\	�S�H-��vˋ��c�#�S��>��|�������6�
��y�A�>�P)��<����k�b Տ1o�b�㤯���w���[,�vC�r#!����g"�f�O�@�~O��T�PU��Jww���� R""-��;DZ:�I�N��.���\J�޹����7o�aƙ}ώ�Yk}>kﳏ�ėOh����|~d�����f��n�5V��H|U���:^}������T�N� AU�c�2u���ڃ���;��r�q�ym��Ҡ�2�XSp>�9�S�z<��Ip��7|�y����I$ؑ�����T��K@���*���'���@i.Ћ��7�!���7̑}�H���2���3S>'*H�����{7�Q���:o��?���]�v?��qG�`; ��R|�=��Rՙ�����(���Q�3�쒃CB§j�'�^r�`����D+S���_A��iǳr��������~�{��D}:l�;�$�U4?T��9���g��8���GS� ��_��HU���r��0Z���_���� �fj��2[$��{� ��3��T����q�D�즐*[dIˀ����)%��ˣ?Ƅ^Χ�j6�A! ��x���h���҈Pv���Խz;�a�1A����aHx�:B�U}|��^95	��f���D�K�	0S�+��!l�m��N�3t�5�����%�&�^�=�TϖJ���ֻ�仙��<�i6��ϝ�k��Ó�ێ������9w�o��}'-m�5�j�&UƁ@��w�R��e4 	�D��Z݆<u���FO�zVUc#��`0py���F�X������d�Y��­�c�؎��ˊR� x6�-��' X@���v��7C��Re�_��z����;�;����s'�������/7�ޱ9��lC@�]�RlkG}�{�0BO�{�,����cS��^Q�n��*1d�\�@�t�:k|��%Qb>M���T;��]]�U�8Ó��F�����	@�R8���o?�!��c�K�K��7b�ϻ�|h
���-t�j��5�]|2��әv���q�W�z���);�3���"��ɺ�^Y"��oR=�X���4�*�๛����B��S|}��DjE�	jc<��x>S���x��&g���ȢFX�<��V�c�_�)�ٟeEg{�_��2���ª��v΢m���������]eT�ѡR��ҙ��b���~�����~���P���x�F���7���/	���'��2���'��4h����{����&�lx���	xj��$,^�Q+rH��䕼[G��Ʒ�mj�@�dq�*���j5����2��'���}�nw� D];�L�|f�'�����C{��_9�ѯ�0B]s=�Sqy"l��e��ne��CՇ╍�2�� D�
u	^���^�wa~��x�K7����ʔz5��ڮ����-�v��DۑJ������U�tzl�Z��#jp̃<�q5n76`Y"#X��&��0��4�,#:�];�uSG��o�������Tq�Dd�rB_�	k�2��? ��(Zm����Zq��8V����3�9�i�gcuR���Zc��X��!gs�Z�]D�7}-F@�Kl����,�u�d��$�ըV&��,���N�.��#�I�{����f``��b��ݕ%*Y����p��[���@A/%��{z��齓�$i�lG3�e*��u+Cm�5�Z�P8��ǭ���{CÆ�]�֝K�������Ʊ�蓗63&�p�r��53����<�9�F�,#*̓�-3/�b��9�lk6i��|/��Z�":��ya�Xe
�j"Rr\�95"|�����94��M�(�Ff�u�\�鋞�SxB���y��+��_��R[]O�|�KG�BVե�E�&���>�l)��ky��@�ы�(� )3���H��U95�Od�=�`:s�R���m�
�ra?:�X�E~�~��P#��K~��iw������'Kچ��Y��=�S���U�����>�� }�m%�2j��rNo�eH�����F�*��`���:�	

� O���Z:�b?�ɒ�^A����x�h��K�;:���~!���^�GM�}��J��a�2���ճ?�\�J��N�k�a�~��1�R G�ݎ�&�j[[�R�F �묅�KeX�J/9�vV���жX��/Pqw�iA@�ju9Ȍz/���o��'�NX)��p���!�.}�艹�BiT�uT�Z����Ͳ�	,��A�gm�z��>"zU�Jbve^n/L�<�qp"��l��s-v<��kR�p��i#��j�H(��E�Y8z(A:�8�����Y  ���� A�Z����n+���3� �S�]�qy��]�qΈt��B#ʿ��<�rct��F������v]�&��XZ�ř�ńҜ]5j�F]=��"�$�����L�ղܱw8s)uu��h��eCl{��b�\�!�L����_�r��\�����b��Ƽ����]b��>hke�~�?0]�<ZE��-�?��ogT$�b��aa�n/��K��@���{�C���������vZ�ŴuB:�|�\BHw>v�UR�c8h����Ng��fcپ����N�T>A�b_H|Vqm�@ާ��و��}ҋ��jܠB�k�s�"��c��+.HD�q�9�6r~ ��p��I�16����o�1�X
� �6�ٝ�g	��d� �}|�����4������xM ���~Ů1`3HapT(�S1j���k}^ݦ��VW��DJ�=io
7onh��'2��-l[�t�1֛��5<�ڈ�*� �$:ڝ ��ޫ�]ڊ�ր��3J�̴^�Ӿ�4�����^�����gw�J�`���J�KG�J��V3���@��+����u�f��d�E�mlN�G/�9aH���>y2C澂?b��K�xe� $�[L�+O�э��~Dc4D�WG�0odx��.J�0�	�O� �[% ?P��߀��P�a\�_���*S����w��o]c 8�c-�M����0���'e��1tz����J��㩖�|�H.�V�7癩`���e�-��/�H#&L]����|pO�3���|����8��Ԉv	�㟌�}��F5��/Qs�=5ט� ���� M�a2%�˃S��8����n�E���̽�w�!�*��'$f;#���c�Ly�=��YQ9͸��5�}
�|2G���$���=�=���k^�p�wZ��_���hX����b���;����b�x��Y���3��@��'�j�~���0�(i ��;�Ѷ[Yd�d����c�ei3������PyB�"|[~��Id^ �F>}(|��~F�6)�M�k ��c��3�h}�w�cs�p����k�R\�:U�b�/�O!#�W;�F�5�fZ�m�U�ʮ %��;�.��?1Cb���� V�Đ�v�]��.�˱	x[��pc�Y+x>f��M�అ $ ���`)���W5����a�$.��M�^��H��4���7vx�Tr`ч�y��j!|�v:k�v�R'��^��NED�1d(�����w�}��]��C&���,���`�5�[#?�Ɂ�3�0BQ��zx�����a#/��,�1� �d�w�g�P!��pK����A[�ʳ-������G2�L@GdTN�$Ⱆ��0a�m~/�#�0����,m	ދ�D�l�s�n�$[D\�>̋��o��w�t���e���5�ց���?t}L�%D��9�v�L@8۟$s�;aD�tԹ^�ę�Փ�M�p.�>�T�d��\f�&pTV��F��+�lR���M:�8�S��} f*��#ry��ϓ�yL�N%Ӈ����x�H��# ?�6�
�}ؓٛ8����`FI(�-Wޮ�}4�7䏃@�1�h�W��5�r�F� :�#���2��I�2����t�ƍB���eg�����m���^�v�����k����#�o��͗��g�mU���'��)�]�
�K���7%��I��5���a8�,90@��΄�Iʽ��\��fߩ����Z������~���M�MJ"q�	}��0i�W����8�1$���
0�4��rE��0l$w��3ev���۲�����v����0�芾�S�ޘ��9Ğm�F��PYEd.S��8�`�%����z)m��Ƃ�/��x~:M4�)ݕu��a�����p�z)+@�&���V�]�ۯo�9���3:�-+�	s6{�l�O��Xz�$�#��Pv�vU�G�KY��}����;/N�mi� �y['���{|��D5$�{.�
K�k)�1]��,����-!T$���0�X3P("������h}�5*V�J�i���{+:��/FSPdJi{;)C'|�y����F��Q���ꄍȢ��$HF���y�|�A���Qc��B�hM>�Q�"ڵ
�����P�����	�
s. �4t�!�����,����~��3�?���
�'u&��{��9�����7��qMed����1��S���Wl�k;� �R����<��D^^���* ̔����-/�).�X�����f5�.V��wi����Xچ�/��x�b�yŠ|]����pq.PQ�5��i ��1�L�ͅ�>g�n�Ã��uf4� =�F_��{Z��6��$�u��*�;v{��}��Ӽ��7��z���bԺ>~�2J��x��m���%x�����2Vl-����yA��c�7փ޹KQ	�A��D>��9�S��T)4�DJx�2#6UKn)��	6
���z�WБ'��v�l�?pI�Գ���*�;���減=KTJ�?�����gӔ*��R���6�y��6�U��C�u�����jG��P5si��i;�1���.
����)F��zx����bZ�Tnq@0�aw�\��2��!e�!�v�SL
��."8>^ӷ��=e²քgO��vc$���!���'���##u���Cy����+(�_<��=�e��@Ν�x�BTG�T\�̣�b�g^�䜁����L!�&���p�Uj�#ut�3GL�kNŌy �G��^�GC���:��,IF�X�g����[���c^8<�/%�M)�Qq^��w�`؈����\��SV�r�;nøߛ_p(W�yF���Y��m����S���(̍b�ďQ��vk���� -��݋�w������qF޷�,RCk~Շ����El:�|�\5Lt��cc)|�mh��T(��,��$�ܵ�ˇ;g��� �M�{Peѕ� Hdj��+@x�p
(�$�nQq��!ŎQO�UFLǿ�V�彖}+��bwIde.�'t!�p�l�ܹ�=RSs߆�C�~��{Lr���f!V��87)��64�UWd	C�~T~eҊ��'#���^=������=�!���/�g���U��F#�X!b�������h���K,��de�}�ȯ�.n���D>�Z�9�a;�ZSĆ�A0 �V/��R{��x�R��[��y�.#G#1Ֆ&��e��UU�})����֥*�4���٦�F�d[^��s��
�ҋ�傇&�?pT��(T;:�K���Ө���H�E XF�v4@6����㗗��F���s#q���d��P����=J�by/͌p��]B�¦�����t��1��^�7 ['�^4a@���/��,�Ml��/T��ܯ��-�"���n�&Z��&%��%^v�F��(��b�g�V�d�w�zO�W\r8��������S��}1ެ�A��F0����>[�G��dZ]����Z4伣U���f$���ejn���	uNcQ���ώ]k���E�xJ����*��\
A�/�5�@n��fbُO�{����Ǿ3Ŝ:���1����M.�,���� ��o��k{�n
��sT8�]�ۧ�]�}[߬�F+���hU�`\|-����`ťSo|��T����`n�3E�l�+��\F�����T��˵��>=�Vibm͸X؋H�+5	���| n��A�V��~�ؓμ�x�`.�5@���� �4�*����9tHJ#O�`��7����̚bқ�J}��'�mvb�Tk\�B_����T(1��͚��o�~�,L_: "���}~Z�9ѣ��V��d�����G�� �wBM_W��8�!���.ms��&7���?T+�?��}]�,FǙ4�D�;��ͫs&��_=���By-��m\��c�x`ol��8C��I�s�u�X�C�o�^D�^�5�P0�����z��)C*�eJ�P�͊Z���N�S��DC7�����f烺�U�V�{L�h"dp�����(������YV;xŎ}�I��y�:k�<F���8bް��0�0]9R�+�-��<����8Q{��O'I��hۯ,��	�!�E��^^�nJ�T]V�ϛ���_������=�|��6����jVbV��%��BJOr��D�	��K��>�E�?�{�.(x����ח� �i��ڐt�|
��e�GE�d�sy�\��;� ��)Nq�?��N�����ܞ7�����0J�?<^g3�l1�ҝ]�x��48OV���^+���<��wtT�N�� ����qF	��� ?�%_��˂BG9��:\i�~(�~�ݳZiq�ʧ>�NHZ���hqGE�R�N0GiQ#}Ztc��H��Ώ\A���sԁUF�|�(]GE�/n�ߙ��4����0i�����ƧXgK�d���d��w�bU�)���]y����B�q�ʢ衭�_�q�'���`l@c��b31l\ӕ>+���G펉�O�&�6zx��r�����:ݒNj��w���8ۻ���]�����f��ӔF�OR՛;oE`(�J#To�����|,խ��#�d_�~<|���/K����Ե��1��ݔ�n���6}�ߪ�)�C�oC��te�$�V�&�]P��7}���¼9�!����Z*\ p��y,��
�uWam�6��4iPG�lZ���pسu9��ލw�Tqm�d��g(��U�q����^N�:���q���o�����j�@=^����d�������ݢ��ߌ� f��ߎA�d;���Y>���ڐ9���V2��@�@N�tD��d|.����HJ�CG�������[��[t��݄ Ճ ㅓE/�c�yZV8|��9#i�?��Ҍm_����k���J��( P����.��W�~����Ɇ��<;��nd6�P��6�V6�T�~~�D���'c`��}��{�M�
Z�t�,��o����_�*xiu�ұ�B��{-q}�E�ߦ����D+a@�HJ�]�����޼CO�mYt�4~C���7���A%�y��5	ߪ�Щm,�`���۟񷟌\���󥮙�������Kg�}��6�,���O�R�3ʮS�K�Z�N��1
xG<7����a��4c1Cm�@�rm���yG县�Z��j��K���/��%�˳�`A`���v���<Ðfo@�����̿Ώ��TF����8�*n9G�c#�1OP?��F)��&s+O+I5.���
[������t�JfU��n};��m�$��������V2�j*�{��Uk@rw6C���1 "�rKI�,�l��u����a&���m�	���O_n�2����?Ո<���ӗX��[x�6l�M�C�|��K�V�-�;�V�}s��W�䐅�,4 g�������kq�k�8�c��8l�L_��5��$�K�Z���ɿ����bU��[���.����ꘐk�d=�eM|��s1Dd��+����>���O/�%�c��)�o�� �t����s=�:�����-D���׳9��]Y�P�c?��9`S����)�*���)���-��ݨ�+����rӇ��¼�PG�#�c����w�^����ڥ����{�l�ը)~Ȋ��(b�	 ��/K��9���0���ɭ=?�����s��Շ�1��?��)6¨ٙ6�/3-�d��w��y��^ 'Ӱ��x�������� ���nE���ƀ�U��a����P�|�?PK~��R){;��0ds�����B ��P%�4_�N��.}�Z��gg� �a+�5�	v�u+^z]�A�W�@p�9��-�i�oƺ��H~y�z3=R&P�[�kW�T�(U�q�6-[���]xy��1!. �R�����'��j��> �;y'%ޡ��L���
�#���v�����^�x>�[NW�x�d$h��� �����_ڛ��mժ
Ŵ�E�Z�9������j�Ƕ�^�ӛx�\�)Mn@h*3��b""-~ﳚ9�F�'����״��|�W�j�*�#{�o?}o�� �~Zl�e��"����`1�Jq�	!�
 �J,�#6���P�lBب�[���w��|�-�J/5�Ũ� k#ޚ�g�Sm�jz_���S����t�F���ȯ���1�|��}�}3�.�T���P|�DN�-�9���ˈ�g9��F+�n��p��^�����S�ÁP ��jk��#F~ ��S�鴗�m-�WQ�	���τ�G�isg-Y�+2���R�~'����i��-��q\4�&h'cyc{��N�~�V��4��ۏ�[�e�"Wü�{BQQ�v�Јx��Q|��G�!�Z+�EE�'|�� �넙��ϘSF��t��ÿ�g���k���02�Lavj6�ޛ%:ig����)������^w�dę� ��L��;ho����+	�yPh>GS�[�b@�i�%���������AT/>�}��2�/���#���*�f�ax�FR�l�y�����}i>R|��>t���t�̳:��?�81N�Kf��ݱ��4L�&� ?:�5t�Q�>W@r5�BM���h��S��'�['�b�;h䅆툔a����KzeU�̭�_��D9$5*��u��N�3��nL]!���f-j?�ɄY!�^�t�=����!x��~��N�i���hb�a�r�Ɔ�[B�qN������&#��>C��X ,��,��''ʟ<��I��\���������߁�X�:u�Dr[9�x��8���O���~��T��G��g��E��Q� ?׫�%)�4t��&,��J_�t�lEj�����i�9�3޶�¶��� ���Wk��|��6��'O�+�$�`�\%��� �:���4�1�(3��*%�`6i�V���8+�ѾK=�y=%�4i�iy��tRf�"2OK���ĳu%E�^��7.�����*�OV.z_�+�c�jH	��J�+����$�ȅ�m�_>C��m)�I!QU�eg.=����Vh�ݿ_�2�
X�%½"�b%�P�1�?���^��/>��4o'-k�{0����:��J7��"��n��p��,.�Ҿp:�&��*uC��Գiw>Џ�h�h'��T�d�Yc"�����QA�s!<�a��u��(�U�`�`»W��D��}:;{�1�J�5R�Q�I�c��TR�4���A�o������o�� ��lB�����x���f8^�M��r�g
2�Lܭ����LM�|?�.�g�@-{�qsb�1��u3�%zvZ">���t����SAW�'���n?ݚE_y,��)���g�x���^R�Y>�����}���b�W���%Q"7�������V�V�{�MT�#eE���:��ր����o�ς�d�=��ۜ+�ѻ�Ab/>��nJ��}z��75 ��}��ِy�x˂�Bqs����?K!1�|��>��б�`��2��$+��(ʧ/��Dk��
�gT��K��ZX���W[�Ic�ϯ/'ť�!�g*������7i��Z��:��@��r\�������*�'>,$�+\�c%�]��鑖a�qT�8{��U�����FY��$�f�$cf��BM^�u��r��B.�}�`UO��E\�<������%� l*��eT��{�/�U.�Iх./�l�[g1���w�6�t/���i��ͽ�q |����=P��=M�s�Z����t8!V�kW=��9}x;ΰ����E�4 =�G)��6`,�T'�9BS��5�x:�(s��oZ-�/R��f=�	����m�:��O��N,'֦����g[�K6ۘp�{g����XU�L��R4GF�	߫�_��&��:���+�d�K�o�~�ه�5|뉺����8�v<�4%1K��-���;a��f(=ᑑn(_r݋����/��})�w�d�J�y�k���^xgIMɪuKx��+8����Bʏ1Q�#�$#��6���O�L�����������ܧ�\��G���$�E��k2�?���Me�/8�����<hb��=�T4���Xs0�X���s}��zF;��]�Ӌx��1Uɏ�y�Ό�$�/��w]Mf����Yo�"�X`�}��-5�i��"w[��z�X�	x!���d�Y�<�i��e;�l/x�38���/9q�qS�y�7_���X7�S���qx���(n�������剎����ⷉ'��;���lns�����]/�DI1���ҍT��	�o
YI��c�؀�����=����1���*�������t�v�[���3X'?���OlJ���2Aj��e��ߗR���Ս瓕"�y T�T�@搸KgBY�qr36�<M�)��(Wå�ޓg�:�	��RY8�ת�jd�G-L��w5��d{�WS���Vd�v{���a'<	�#�Ș ���]Z	����~ъܐ�n�Wl���m[�;�4>�b����;j�6�{r�?��o��|=�<\�ߵ������~T�0Y�"�>��J~���RX���f���| �����[j�S�`k��ݝ&c�s�֜�eIi��_mv���9rrWW�9^p���?�,!����y��
A���e)�-��5)���zn���<�����Ԇ2����f�p�3G���1}�Ḋ���7���j�i�g��~H�C^ 5���[BCml�2��t��[z"���T�ۄ_lH���B��rG���.��)��3��S&Q���<��X�!���=C������je�4	�ׯ�=i����w,D�bX���8�bO��\�^��c�Hq�>�b��l���g���Y�6����Q	`��k������D+97/H۩֟�|#�=��G�yҳ��� kǊ羬�3럆��ʁ�M����i��1���%���&$^��<�^��N����݋����b�G%>�ֶ�{BC�e`��Q;%��p&�4F�h��"]M�9�sw��˦ ���C1�
K���I��ι��ߍ�{��N���5kQ�n�)�<Լ�ќ��Dr75F!CU��_����e�y˩�B#n��� u]T�yo�]Ђ'gF̴�ia�S���]����vY�h�V�.O��z{�g�;{Ӫr���h䷺	sXZ#q��p=_V�כK����&�Gf`����t��"+�9�U����=�ѵtρ��.������=�Y]vn����Ã��L;�f�p�ڋ����d��p�x?�x��~��R���R�t��'�N�r"�rF������2Y�֮�@�)���[�E���K����ZF�U���Ɇ�A�&��Bg�n�H�wFv�7��߸6,���1th����~��蝶TEe6����t��i}�W��l6��mq/�C/��G F� N#�gq�"'���8>_K�d����WSW�C�P��������fF_�������X�k��B/?�ԇl�IL��D&�۪ %���#{�.s��xN�Lt��N��F�0硙zD"eN��C\O�e�߁�Y�^O�����zlXLW~���h>�R��� ͩ��Ҧ��~��0�/�`X7C
���4C��w�z�*fV��ۅ���N&��L����^�sS�1�z?�T�H'C������	��߇��f��&�H0�9`GK:sz��2���8OtYg�0*{�
�1U^u��	�|��Z�Qx������Q�W����ێp��>q���ɶ�RI�Cӝ\����4x���6um������d"�9ݴ,��r1]��Rq�䥍�@W�A���DJ=,���V%][M��-~���s���S��͛���lrXuha�$�eӹDrъh
��d�T��&��c���������>6�bO�����0mqw�vI�ۍ_5T.���j̿��Hu��k{!���s�����xM�������R'ݫ	��G�d�u��7F��2!R��Cp��p��H��ﳇ�;��$g�4n��l{�-OO�l���y9���=hZe�=��r`�SK5X�o&ؔ��&� ԨԼ�M����(��%���!B��_�cJMˆh�Z��u�����!WB��� ��櫦�2P�_N7�����N</��a������n�%��pB��_|p�U�,���A�w͖�o�֗fi{c�MW�Y�}�?�&]�);ILrY>q��D�O0�`�R$�iG_��lT�A��*�(��M�Y�\נ�G���.���%��B©��������� �H�7:{�.	1��߇��LoF��ө���az¡��~�<��U���O{����uyK��W����.A5��"��>[M�y1�\j��s3����]���7��@�_gZ�	Pp�0T�ŏ6M����R���%�ԍ���C~�]=\�bE<�n����b���3�;[�RT��_�^���� �h�CB�p�ۭ�F�s���n�C�!gI�1�r���d���څVV�M���"j6�����3�9ƹj|����Asߡy��Bƾ®,�T.� � ���t���2���!2����sq�4Av���]b�9B����:Ȣ{2�i9� �Y�M�k򞳪�H���Y_>�w��7���-��*�5�0^��u����Bm�����W'�mAFM�����$���U�i�߭]}*���Ma@ �SӵM�/�~ь��e�f��%I(���b�m2�)cdf���<�y���l��I��z�򈼓�9���0G�a�f뉄��L��(����+9?�M�^Y���oԎ\�������oGE.�q��N�e���7y2SP�J��Ƙ��H��X�!�åVl�0��_����Dr\�����e����f�D�TAq����E�Q�,��֯��c6�j���'Л<ŀ�g G�p1�Ck�qn=n���7�;��Ȗ���wGY�8ν��+��MI�/:@;mT!o�~7�p��y������r��Λ�4mfՠ�=^�%��� Ö�;�,���SY��$od5\+06�3�����x���n��<�')�u���ߞ�:8L���ֻ@k�/��idx��b�	�m�L8�k�8�+�r�X7�^�e��קu^�/�Ϭ��L����m~طoگf��@Ĩ�ˡ�92�����nV�],Ԩ%�:�>��4 ;��q��XY7'�H&�8�_�F������37�^vȜ=�Ĺ�����g���L�Z��QY:���k�����j��\E{56A���7 �xy�L�޽�w�phrҮe���2!B&�e�J�>�h�^��)<E�(�\�̌��f3��vl䪑��T��^�V{���
fD��#\����矬��i *��5=�k{�'��P�vt��(�07�s/��ohM�u�a���7c�׹�{�ɼ�m�V�9�ҽ��aasA���P��m�QM�0O:se ��*�8�2�RQ˩Ċ.a�|�ɆD���g�Z�q�4fæ��g?�C��e�J�� �Е7cr�f��re�7�,�|.����[�����r)U�V}FM�6_�����ڬ	��Q�f�HD+�⥝#/�'���E�f���D?��	�n�T�|n��d�Z�{{�JW��|��ɔ�Z�o�"����F2��۶�g�՘|W[�����c9P�'f�,"�TCE��B��k�Ä���޿����G16�`�"z�^�Ʌ^;�s����a��#D��0�p��Lv��FEg�Xޕ>��F*G`���G�{3�b�A��)�GX�xc�V�*L0p�7j�||46������e����^ �N�1r��ڐL�v�æ&UPN&�J��+⧣߶��2]���Z�#�V�aD�ˀ��o��M{)�4{s'�Z��%w�<�5�Q��筼i#wu�y��>��y6�W�������/�J%�/O��*kj8惠B����`졃
Y�l��d as�� �B蔚_���&1����|�$ �X� C͘��w 6i��i^`�ֱ-`Ji��sv�8Ȁ|['��(�?��;��zqd���H������/fI�2k/��ɷk��M^qF��o�ԡ'J6_��b�������9x�n�c��ww�֤i�'��:[&�x��ѭ祫0-��T�&��@�B�f�y!�ż���ژ-m�nA��>7���D���e��e���c�x�7�؀H��$W�$fpI��*��s!uPc�̢�m�j�J/���e*�������@0�ԻC����`!����D�?�-a���Zhs5=�O�O����[��4)zRDF6\��hi�ϝ��R�У��ce��cIQM)��M�`ϭ�Z|zd�,�J8�Lw��F������@ ׀ڴ�Er�ٛ�Ph�A5VԶ�z�A
bk�O><�M�\����^��8�;W�K^���1�v ��U�v���J/�oze>^�ķҵ�?k�Io��-w�Y՟7�o�����XX���ɝ�i�[�V�ɫ
6������s-���4r�b$~�:;\�MEK'"�3�j?3��3+��|2%��/w�8�C(�#L�I8o�s-�}f2�z��1=UI��n�:T�8�OÉ~�M��]���%�\�^y�����8��\|@$`�<{."/����V�do#J!�����M�^u#AÖ ��$���݁O=���,T��Y��dK�1�� �0yS����0�yG�Iמ���[��J\��+�4*�L���e;["���(��ڣ�W?J�	�\�Q2k�Tp����q�szH�y�����0�߱iHy.��Wt�t�<L����De`j��s����a6�G9f"7��L�v<n���y�Bڛ�8E�M���'�~UD����b��!Z��Ն��ո_ݛ�\�#P�7�)��'}�el_2�.q.3����e�=����&ᖑ��"y!���#ݔ�oֳ�VH��v�[�f^���Ӯ���Z@0s8]x�d�I2-�u��I�&�����:]�w�G�x�4�`f#��*�[X5�ϝ*�w �}�w�1���'���!�E���y�����T���Ų~�q*l0%�.�pŗA�ւyE!��l�w��WV𩬐�k����l�)F&�9�7����r��LUU��,3t��N��);zp�	&��*(�,U`��!i�����Y`z�1�0��6�p%Dp�|葭e�k8�zS�F�=d�%���Q�,��I�BV�2��M����i2���M��18\3�����=��vL�.R���̪�h
�"OHG�6@0� .��s��=~�A���{_"#oS�ҡ?����ʨ�}O$��4)��r�+ U,�rNcD�W���+�*��ӡ�{�;��;�-�=��8�yW�)�.�/'y�u)����_ג4�2��	=,�͡v+���	�ٛq���3��	oq�[RB�&l�U���#o��Rt\�v9�0yޭ<��`�@d�����ͦ�8x b�����k ��D��r� �)Ò%t6���l}�����ߢ�����a�B���
��=G"r�Qv/rɄ�?�T�-���Ba�%mi�k`�i.�9�wv�z^�h�F���(L,6Ȼ��:���D�Q^9c9�x6	t+��v�ʉ�W��:�!/)��K����F6�*W؇ �+�������q�F��Eڡ�.����k?�<�_��+����h��"ϧ�"!�J�,C.(���νD��0��c>،qؓg4�ڣ�`�D*Jl���#uue�(~��4��N�~<�fz�'�N������冴GgQ)��Y���H�^��]A���@����Z�s2����:�����\�t,�˟Pu�ZFudSP�6�3�X`����b��z��g|�( >�ߠ�p�S熟�i�a�
ı�ך��i}�/͉?�R��j n��BK��|މ�K��2�M7~�G�Gy��;>6y9�!N���+��q��&��jp��7'@i��@�Ázr<Sfv/'��qV����=�D�R��E�}p�f�:�!��z-$�E	ZK��<-�9ij[�j�~�]Y#��m/�mZ����
{�%%S,��:�O"�O�d�r<aNWf��.ۻw1����TQ���"e�����gl%��3[eݢИ����K�	V�T��r%��I7ݖ7&��Pj_�3|:�rKF�N6��w������ W�XؓQ��{Ew��L"5�W�����4��*�/���:���ڙ>"5`�+��:u�k$-G	S���sn���	a�>:G�;�� ��U���3�$V�I,ꈐ��`�|��-�A5�a��Y� ���!���1[	��3����Kbj8H>	��cU�a�;m��h���aD��]x��4/67�VH\�3R� vC��Y���2���k��uC��Ϥi�.�j�٪��-���{��U
�HW̯s?T���L���z���<ٝ~�^?����T3���F��H��?x�n��#��Lm��mx#���1R���:�f��%\oQ)��JlƝ�7l�,*)�_弊*��3 ���z�:p��������{�o�P�q%(�/�P��Ҡ�dr7gB��\'oZդ�\<�c�z0S8]loA��W���T�N}��o-�^Y���[�ã�^�5	2�3ZC}���}�����.�	9�Jչ��Dze���A٢�Z<7
��_�R�ϐ�v��B-\���QVvL̽)�-���$D	D�,�`��U尘gi�$��
L���_`�,��
'�x�2�di�e�������46u/���N6s] ]_�HU?�	L���<7�{%���d��?���4�:5j������q�^r"�KN��PAݤC*�Z&_l��9���%K���x� RR � d+r��s�+��T"�m|����׃r�B$>���B�J{?�f��9��f��k�([p�#j�'��7�)P�q�޴� I,F B6��ex�����F8��13��פ�\��]����U@E�>��[@Ji�nP��.��A��D����\�c�󻋿�w�G<���y�y�y�wGر�݋�_�?���Y;���`I�T��=��#�����6[�>�yhv{Ȼ2�5��G �5���5˪�'�+��-C\�`iI}�	�i�z�7[uA�t,���D�Ju!���ъ�������H�yҒ��t��*?��:@[ =\Z �j1��0�n�}vӜ3����_�qcoBlR�!{�QaE����E�j��=\D���~G�aP[{���Ta�:~ܲ=�Wf�ӳ�5?Q��2URW+X^TJP�"��p;7Py��YQK]���n�$z��G>bu�h�ۉ�E� q��@�����N�n����֏4�ی��
�*])Ӟ
�Fi����v}z�Q�}y������)Sn7WVS�_��ō?k&�ҋ"t�ݨ�M�p80�X��$L�O��A�_õ�P�R)a�1�ʛ���9�&��D����'o�"@}zN<��[����֞�-�~?�]D�����B�{���?X��{v|.-4���hnX���X��_��]
^������Vc���G͖��󚚤9]�c���Ρ�$ߞ��8؍�.�m�Is	���t��s�V��s���cd�,̗�rG���.q~ b���ym)�υ�I+Hq�������ϸ�H&�fj�ʐ��
��I��ɀ+�^��;�*���D`S��1�ƥ�N�G�r0���A ���Ŧc���H�Q�4]$�џ丟�s[��m7
)6
=(���u}]n���S�oI�(����Ȩ���.OR��׳N:pձAg��CdoE���eͻ�YR�S��u�b5�ߴ;����NM�����U"����`O3�:�m�x���#�Ys��c��VM��`�|���.7z!#;��̤ǂ�׈�������Y
�l9�����N?�5k �%��(l68K��P~�&s�Q�3�&PP%T`�`��f��T��U�cI���Qb" kf���LSe��W����E$������o�Tv2������n�'�;~B�6�M���%�Ǖ�;z����ܹs��6�A�`��C��)��>`���=�}���Tι�}�D��qB#��ۼ'Z>��F.^a�:2P�V��ݑJ��W�s�^{c�d7�&�+%l�{�"��z-MLd#9+�P1���"G��)��>����J���7/?��@r"�q��f�T6q3�ݳ֔_���p�*�Ň�>�?l�W��۠���Rއ܅Z<\ ��' }>3��}��[�D�5U+��kQ~��f�J��d��WA��`�[�.��`O0�	��j�j�g��s��)�y(o@L�*Zw���E����,�Tgu~���
ے�1߹��&�N�-ov���f��\��"G��nSC,�ր��ki��>��I���3����'�H���X ��f1u�;�4����Ŭ���~���a:=��xOB�nN]Y)�d�<�@�Se\Xa��6ﯖ���륏g��	XT�hēK��Pm�Do�ԋJ'B��9�;L���9�SŒ�IL�p!��l��Q�DK���_w�S�G�qػ(w��Ү�����R�_wr�U�S�I
A�ِ��p�RuT>;�
����+����Qˋ�o��M�Ο����=P`9�咷��_r��P�W`ć�E�`��ǫf*��vCr}�/�� ��(�=
b�>�Z�3�zAx9��iw�B��&��s������
u�P�Z5g�l3Ao
"��Ɗ��Q+}d�k���D�5 F:��睳=Rp�|E|'��^ڊ59^aY�d��<��q�����Q?/F9͸�3c;������?���|�n�
ZE�/��o[�(lM�*�n����S�z�Ve�0�ɸ��S/�(|%�WF�;�DS�En��!����V���t�5�ϙ�g=a� 7'�x"c:�&9�m���%~��~Kp�R�*�Sܣ���;%��Z#A�xCe2;���wӡ������5�?w�h��*�ׇ�l;�ۣ����m��{����Z��V۰{�0-����(�%]�g�����ͳR���aPݰ�1�%�w��DT?��.������tY�ٸ�+��]��m���+ʮK�O���6�����J��S�ӘL(������}=)�;#���6C:V4!�"�y��q�K�-�4��ƴ���Q�����?(�{�l�nwtI��&��oj(GS�	*�a2�hհ�HB���-n ;|l��ޱa$A�ئ}�	,Xͨs���b�� ��q�q�(���QoX�<R�wk��o�@�nu�zῸ�~�%�﷌SVS ��km��!���J�1��1�k/�������P�3���[��Q�r ʲv�%�a�R8��7:Ȼ./�c)i�4{�y��W�ʞT��[SU��y�!��g������x��ٟ�:I������"^�?�����M�eP��2�!j{�K%4�lv@�B�[�@o3�J�t;����H.3�;�f��9�~Q_�����k�ť,��L��K�Z�WF��Z��b8�l17#$�R��/'���y�a !L��w�eCQv���Y ��O���T��Wx��y�u�����y,��L� S7_YJw�ByH�캖��Q���nMY�N�/�%��T�xo�ɑ���O�h�d_e����_�$ ]���=OΊ:�m&�`����&!���vY��� �#��'���S*<az�w�J���^���Җ ��T��H�Ӝ�3�_I�'<�P�[����a����O4�!��Fm`���K
\��R�3���n�^zR�&K���|��+媎c�2���
Ȟ�j��khI:�1��rT�5E�>h�u�v����|]��JMp��ν$�����������\
�*(?5{)&Me� �[�w�	΄�5��:x��������U�I��ن�hק�1�Vm��57�Ⱦ���d�[�m�?��*Nϩ��W(L�
�� 
�$���Eb�4o&�\�^���f;w���nӁ�7s�I�l ��5�����zQں"��5jX}zݫ�K�����at��T�=޵y������������m�*c˼�Y���^�rWwDo�M��`��T�k�l���ˋ{�a�
nam��u�WX�.r��5;�8�.fgD���.�A��� �̈́����	5��FO4 �X}I-����D`v@��x6S<mVw_��ց=�#�B �̓[@a�H��D�j��,;G��!�DWhY%���2�D��C)KV�����QX��Ϡ�{�6M�#ЪS�r#}�5e�]���̳�>��\PIg��q�w�������%�#@Ȅ&1��K6���fyw�< j�#R4�MwE{���;+y|0��0��U���d�R`B{̸5X�/W�x�4s�!�ީ�1�Wr����	?uȚ�C���]�A����;y��x�Æ光��΋���w Cb��uM;��0�컮�\P����#��̥|�r���I�,�M����op�6u矡���Ԝ)��+h.��/���l �w�g���s�H%� ��p�S�>��2�������h�m����I��`j�a�qo����O�y6�I
���ￅ\����rh �&mo���m[˴��:��D�TPc]�fu�]��&7����$s4~H��� �3�x����b��Y|�d��0�ZB������$s��j��]��ؽ@��
W���`+'� �򛻊_Y(	��D�2]��*f��t����Ӗ��ߧ�cM�~���Tɯ�Ca�X�R���r^3ﭫ>�2e����*GU=���t�++�v�_������Q�ռ�Ű�ϏА�W�Kf4mh�Sm��kD�/��,7>=�6�s]�q��
���TS��Ǟ�ŉ��|�T4A�̊7�F����������-�4�}�<��V�}���{%ۨ����wŗ�ַ_~{��䈠���o~�s�+�]���Ex��jx�'9Ǭ��u�9E�#K h2�D}!J���G.ʋ�#/Z,�H�g��6��o��x�M��$f'�P_�'y�ߏ��?f��)g�/V�v��qw@i��dqϪ��ßZ,�&�t;�]w�sG��[c?������,��㖾N&(�+��iv]��S���,"� ����yt�T��5+q�0�ǭ��0�<���w��_|�G��y����|�e�@�x�R�5��a�b���J���±��=	����	�*4�	���� �į	i���ws��O�$HY󺕅,���p�X��C`C�ZB+>�{pY�²�>E�ڒ�+��/xv0�Ċ
�{[��:�7���r�����SI�O�Sr>=X�s�����}����2xT��$��D��:�U�1jI�������?��EѹI��C`tAO3R:�Y���4����B.��	��@&"��f]��>�ڞ�0��W p�}c��J8�m���C���s����⍇���<�H�?sch�}	V =���`h4�Q�UD[i񓿖���^�r��Dk��Y�/wϧi5W�te�n��)�X��.!2I�UjW~癸f��<�g���hA�CS�l�\�=��i��m�ӟl�{�oG�P�9檁��P,�z��&_n�}�㗴��<-�m��ۂ�D�	�=���������~���T�����6�/�J@?���h7���xƞP:��5�¶V2\�k�_�C�~a������Et�!@�cdUm
�[�<�%��^6[�����lq}�BbA�˿���j�̭G��I$�h0@��g
t�d������M��W7߬-�߳ܵ�aP�pT�k�:}0Ud(m�Աt(�k1���/�������wx�4m	s���x���Ҵ���x(.�
���Rg5D@%�d0%3*a�Vr >B�$ ����h�_�S�s����Y��ᵷ�a�N��U��}��ѩ※�������(tw��#t�aJ�?t�\��d	�{��x�L@o.V��׺��@撮��c����I�L���nh0����^�GD�O���J7fb��,�o��,/�
��b��!��?u+o[�П��*܅�!N��:�0s�B^��$�X�}�s���\�0N#@X�W@�Jy]�r�A[�i����E�Cm�����������Ic�F?��I-ۓf"p�S�0$wg1i�6��/��k.��%	qm�w\J���ҵ��v��yZ��=p�~�k��l�6�le����g�U�n�u����O����A�G?��^'ig�<�g24���~�D��5:��s��Đ��ؙcT��r�����LM۶���fןe4[xHE���N;�j�����B���|�O��'Hw��:R������q\������P�!�<s�ω���-��H+1��=���*7,�A �%�7�/��H|0�]��>�b��Ex_/Â�9�C�r���݁����y�d��9^��8�����O�M#a�r����W�w�T��%�=����Ć"K��zō�l�ڑ�P� =����� #�l�	!\��C�F��)�j�ޖ$Ⱥ��>���=�ј�ܯ_eq%[����f����C�"</s�/c�Yx�]b�^ R��g��*�wl���V
ѓ�<�UET[��aZ��9��:]����$9r�j8ѹ�R�H���Lf���H��$��� ��r�� ~�=����3긕�&^~��F�����M�Y��WЃ��r��6�t3��͚�Vf}TNoO�I���������sq������0=�F����zm�|��z�Ɨ��>Uˆ�١�m�fO�yC��ǰn��4sg�Ƭ�|���eh|5���nA���~����i�u%׷�lAL�����n{�T�*>f����]�D�rG켤~@��o>��z�"J�Z�}{�h��[Wg@��\$�:����5|4�y��Z��i�>[�W�G%�M������CMjؠ+2=l�ea���_���SԨ�[o�>�Q��/���s���_`Ӝ�`.��7�o�����"��s�V�B�F�sx��,a�T�%�L��?�4p��$���o�S�?T�7�g*kq,P_@j��$Ud\�n��gy���㒔Kd�Ȱ���Pae�4�}i��#�Sd�'��%�\�8�����H���t��ڹ)�D�a����vν�����������_���$�������C��ta�
����K$��`����{3e�¹j�N��$d� ���m�(�k��CD�`�E��C|�﷋�s�]���S?A��������-\�Ǭ���ݝ��?B��� O}�	H,�y
q�W������X����9�<9`dvh��{��z��I(��șeok1��	I�pT@�gu�q1$1`��nQ����`�<�H�o�A�z�|�B'��K�ɳ& M�[ض���g|��9 -{2l�/]���}+¸q�P?�}��_������� ��.qi�4v%��w"?�����D�e����,�}��~�^�~6E�)b�?4d�C�g�{T2'
���+|�{�}LV���'葾��!٧�,2��"I��m�P�A���n0_��F�����Ud�.�`���3N��e{q���S@q�j��o�w�o5���g}5C��Sl��ǃ���nV8�G��V��+ءx��T���5�_|�H+o���1A
����F�	Cg�P�씿������ً7`e:"��<������~�ㆥK�($����nΰ+�M�W8B���G�y�J�;u2�~::7�UM����o�vĩ9ˆ�xgdiA�s��q���D����F�	W�FSA�����M��I{���g�Ұe���{���w;�&�IZy��Uv"�Cϡur�9!e�+Ү���ŋI-m9��}^�%'�Yن����ѾSU�p�&��]�)ǵ����Y�|��ma�s�+��b�\�k�)za��R�]N�hP�2�k�r�@(e������a���B��Ǿ��w~NsF���y��*z�-�.��ـ@��ck5y3����̶b����Ә}	��������#��}3]u���ֆ4�w��tSWp��(�ν�*=3q��{�����-��}���h8K��70#p��8����V�m7�6��-9��3&�ʥ��i���>K�Eqh�W�]6��)�x#�hE�Z9IL�^XA^� �n,>X���!���'hW����5��N,��A�c5�����Hd�Tta��/Q�#�3g�J���� �
M2�\c� m}*��֗��i<ô*���I8�@]~V�W躵���캺��Զ�'l󫼨��{���t�����N㋿�Y�Z�xa�fTԜW��/帺�#D@@�!��K���ki�z��F3�-'2ܑ��'r���4�
��'Z�I�<9D����"��l'��!@��u�ր�E5�zi�q��s�k�qȳ����);��B
P���%���z*�7�{<#:9�~Q?��	Fg�å<���xLZQ�
6�qdoU��v4�P���o��	F\TQ_d��Y�_�V�}Q;M^uf��Ӹ������7��;�eq���+���s���G�.,s��ޝ6'����LS�@��kM����R�&�$���ר���@PN>>�%�0��A��,��F� EE�JE�y]��BiM�O�2������G�<ά`�	�����'��?,]�8���t�+��"HoW�pA�Tvj9�}7�x�?-N,ˡU��| �LN���tX@r��R�ɟ��2?S��Xۍ����ͩ�ޔ]�C��p�����Q�A��%���h�G�c���@���3�#������r��)���0��'Q��H<�7䬄}�8w����G�<9��Ǒ<y����`S0��0N;�PT�K��c��A{�#V�HZ�������I)ք;b���� �|b�����d*{��d�B������,=������ۡ�7���<��"A��>��4�my���m��[�˕ \+
�\)Y�ua�- I�q�,?q�M��.�K�j3��������^�f���,�>{���<ܗbı�'l8�5�EEI�ƾ-���$ŗR��Og2WBmWIMM9P~���k;؀o*0{7T�	��H���ǎ���*4�Ȅ�íFв�ܖ�T��z~���k�c[2<��c��b������|6Ԑ�lK�4>�nM�h��:I����^��>-j���v��i�������1����:��دW6c	���L.�k�͔�S=���0Xq�W	:������]t-g[�#Ϲk| ��V�G����}ݛis��W�������׶V"���2��Ϝ��LuQ:�Sr5��)�L6VE�T���#0k�兇X6xh�k ��oO͗%�U��~�jI�'�i���l�<�[��b�rc���9��������w��Ȟ����3:���y[�(�xl�0��+�l:s�]\�� }/���4Jt6�Bƫ
ו����,k��!2߃��F��K��i�m�^�5�&�V�+@�C,k�	�-D�/�����!j�g-�5֨������^tq/CtG�������dH|��Fb�$�"������n�H�J��S ��P�Q����T#����)��T�_��V=M- um=S$���>H(��ê}�|��`|��ā���.ԽC]�&,��A�qM�(g��O5B������[�p�Z�!2��t�����d�������<Ej>����P��4d����6���<�y�ۑ��k}��>ր}w�1;ή��kt�r���c{�*iD���%B�׹!��@l_ΐxo��
��`��j�*rУF�.���o�) }������g#���!a����6E2�*�TL�Q&���(�W��֌��*dof�'���_}�D�ٌ��%�,B�7���h���k#��#7�$K��A}'l�J�R�d�rkY�����~��mZ5td9��rjӷVa'w���+bKi��a��Y+�9\��o7������
���h}ҕ��_���]ݿs���)o{E5�bGF�c&<����=��T�:���rFg��������Y$�=�@��E�K �$ҥ�T�J}u�ܘ亱�O�&=W��ǲ|��d����o5E�\}�/���L]�?�SQy5�^;�\�)lj����+�J�+�%�W��X���R
�t���$��ɤ�/�2E@wNv�z2ֽ	2H��a��IQ!0��wc�DT��Q4b�7jrhp�^1#���V�q ��x��I�tG��E	w<�&Sd�ov.�ayp�jrSyF��@�+dx)�Z�4c��,p�,i�+4a�?�;y����<�?��+xz�BO����l�
�z����MYR g�s����*�7��^�����~���O��c�ޛ��	��	_�0��tP����C���<�g>���#�oy�zrC�?g�\q%�ms;�T�Ga�*�f/_~�S48�e�������o��#�t m>@Nx@/~х E����<����D�m �T�c.ZTE=)h$h�Ĺ,?5ΰ|�a�Zr�{��k�EIG;4��Oʈ�N�B`ʺ}�����Wq���;Ǟ��w�eIf_L�[�ҡl�a�.SJ�d�������\qe����Ѥ��l��2>,w��"]�S���p�T��t��X�F��z\B8��~xbx��7MI~=���2):��=#j�uQv�ڌu�d<?
n!I(������P��j��ɛ�2+_\��~����툝��A\N�]��!�Y�
ƻ���� ���H����-�x����q,ya�(=�Z0�1���[���".�7���wfyzaj��q$t��@��cِ������u��o��� ��s���F�#L��wӵd̪B��W�o�@��{�P�3�� �'��x���䱽rQB{�m[k\��ʜP��4��࡝�V�Ե��X2Zf�1�R�D�!^�
��e�^]VϪ�X����Cy����������q��������D�-�Dh�Hp�Nt5�m3f�(�NGA�@!>�_h(�޹��螎���(�4T���z��G&�+�A�)�sI�܎��yot�*#+ǁ��&�2=���sS)����=�`���'Ǡ��[�_�#΂�hAs�xﾓ��L�o��2�@b啧��<�x*ԓ\D�Q��ȫ���~�T�p
������g���X�����X2H�����͜;�[��l��\�t:F�o�8��M�]K	^g���)#�� 9�����W���г���C�OP��~���Z2A?\N�/�@� )�����#�GX-�{`Sq�[K��K��VK
�Gy*��'V8�������4��*P���� ����xXq��{��%13^,<��)otHo�m����u��/ĪV�ցa?V64����e�	WR?o|b|fs���E��������fd-2� z�9��p�t�[����Rϯ�����h�,s6s�JC��,��=��*����	�i-�3�䮗���=��8L���Oջ ���餑5,�H*��B����y$m��U���^���@aڤ^�휐�(=O����ĭ��Ӌ�ʋ�k�t����*�w��~x�8˙vs�I�x��}��z:Αz��4F�p�8������B��P|����,-�Md�ǐ�c42�>F���8�7L�9�M��Ĥ����1�������/Z>�{��*���	�X��Z-�֗��y�#ky�;����1�)�|U�L%�*
��b�Y.���֫�u� �ͭ�o�����H�W�"�/.����	�oG��R���Dl0��0��t�-���& ����f~����f�z�)>[}�����R$bׅ`�w�y2�l`�M�b�G_��A�g�I<7��n[p��?���[���&�:�6?�~��C����!{��<��G�E�b��Ix��P�������E�?����܂��u'���w˕m��t �dT��w���|�k�|ߚa#�tA:�1�X0�����n�6?��)3$��o��k�`qn%�/�y�&��-�h��y��v�ܲ�c̦O����=�zK�3�t�U� \"ha����P(�"n�H`i�z	?�}Fq����Ф.�����y�����D��љ,V�j2(��u��ԙ��zg.���;�P"�n�ac�5�ܯp�:ŷ|o�V��ai�A2�@�S�V��L��4ih�"z-�M��� \���`�~&�q L'��n"���q,��������l81�NK[�%��Q�0D����p����`����R��w�\�A|)���wԱ���©K���i�լ���مW1�>$u���m*L�������YH�J��&OFs�v&��r��	��8	��)��T�܌�N�&D��	+���{�H�/<��Y�B`���xZ�n�-������;�S@�qy��f��߸{�7ҥ������_�U��ڲ��иm�39P���"[��@%A
�G7�����1�ͮ�ݺ�uW��0 1�?�O��|Y�����V�'��[q�;�|���QZ�t���;��w%��ϝW��$����e�Q�̱��$�Ϩ�������B�𷗖�=V��?�`�<*;����>��.�FK�`��s���o(��~jK�σZ����	���re +S}��UAуn���%� ���ĥN� �(�)�<A! 8�"�q��2���'����Bk���;"���fZO�*��.�LC�Y[����)�>/���r�C�]̆V0�:9��]���d�<��l� ��Q8�j�,��v�f����9��t�^��&�Ʃ���C��V<x*�y Ρ ��;V����Z䞧�W��s�����4���;ɇ�e�&�}Po����~��=�?��7�F��F�� V����@@L��]M�kF ��{2뾸\��o�L�j��f���UM����EKL��ޘ�
A�x�Si��y���9=��B���� ϑ
�e)���Wjj3��(��b��۷`�����
�	j�@'zzz$���wՒKU�'b��(7���N�"�4�L�4�!kj��kM~k�Wo7,ede-�yK�4߮`jR��������`D��lEl�ɶ��m_��Y~�o'�&�$�\���������k����B���M,��J�q�o��u�<��V�_9{�a*��d����3��!�9;�J��wB��\ W>���=+�DC���W����h	l���w��;rBo�C&d�?n�v���g���<͖�5���$�1G�����*�f�������?�"���<[��`�\:���K�Ig�s�Ԅyn����Ț\ �JZi�S'�Z��6d�n�@}��+��]�I�Nc g�+�:T[v':4��EU$����zV �h�2��	�N}�*�U���j'��C�\с��n�h�k�{Pa2O��7u'6��4�K�U�\K��qc���#����CʓFZ��?��O~�������H�o�k,B��ߍ
��D7���p�L�Zx���#��DLxar~9r�\�״cEG�)���bC<�&��ږ��zz¿&�i}��d̎�>_�G�TS��lwm���`��Z�{�[v��?�Fv�|-X}�CwqH�)%������?�:�KD7����K5��]�`�7�����<n�J,(Ŏ�K���g濻�(癩��+<�B*ž��J�#��C��!�5I�'��X�,R���j�K�\�4K�4K9 �.B�h%�7oB$+��F��U���h�㮰��V�� �b�9T�����L�3����Em9���$�&s'ދ(.�o���ȸ��U+��yU[{Z`|b�NR����,AUT�!S��P �1�E3��tOS�7pa:9=I�~5g_�e��&���������`�Ssj��t|��7HЋ����έ��"��Y�k�gV>5��㭕Yj�x�����srg�����F)A�5�W1�������n����:�ඟ2�U�*�g�ݤ��,�]�s������;K���0=���1R�>�+�<﹊��7w'�NN�,8�����`8�R���O@0�[�C���ֳ��K����5��Vh��߈w���ڟ�nw��n�^�S���TV1���;�d@���ݣ&DY2�u���:���Y:����o�����u		L'~�੥�k0�*���
U�Fu���i��R�Ξq>�O�MQ��/L��&!#� p�G�l��r�šs��J�G��b�;��
�wz��|er/%����Dm��y��Y �OSS��.��4������	"�`��8Ա��n�]� g��p�?�4�6�����I:��T���xӥ�&ߪ1�y�"."7@=�B(�N�+�0�ӌi�ge�Ҁ=ȁ�W�k7�����cLT��~\�-����⏈+�k��V�c�,���!�����X�U�$~�_Xj������
5��[�{�c�����Qk7��8����E"8��A1JKBA�s��uwC�M]0����1�%�!e�)���<8���o�\�� @��el���D1+���!���z��F�`y�`Ps�FPas3KQw�̸�f�ݞ���s3.���/� ��vv�Ǧ���L`G�t���m{ĄHT:��df����fk��ؽ��g\�ӗ�1�v�v������q�S\����L�-�Q�p�w�a!���_�����>����J����P�s�F<Q�r�I���xs�:�m��?1
�z�~%������r.�l�����3��-w��K74�Kҫv$ȹ+�
ͯ�h��Ĉ��CЪ��)��(���h%V%k'M�4	���������<L,O}W��,�r���ܗ�j ���7d��w
��N���
�6���$�7�A i�w#7f�`��K!A߇��f��~�דXW}u����d_�������S�x,ȵA�V=��F�W��^f��]r���$�r�KMx�2��𕧬�t+]'hȶ���m.�r�`���.M�kN=c.B'������`p	9����P�J��%"e�<��J�R6��%TS�h�Lp�f%�����dH�z�=	:e���Q����eY���{�/]�S���K��V��~�';��~}��LCA���$���t/ދ<EdDCN aG
um������Xj�`����Oa�� �ʈ�^��B����W��f� �b*l�O
&������_D��q���N����Q8� a����)(��C
�7%`s^g:��@�?�c*��2韃�<L�&��AV��(���i0s:�^�-��ľ`��!���]�8���V�6�� t˾�%��sAO�Ȳ�f?t~��_j��<��D�9���Q=�JG@	��tr�2�c��w:7��p�觰�G�"xxf�m~`��L�{����)��PM�?S����?5xj�$���{ء?�p	R}_�v�<~�9��c��/�])0�d[�^��_���P�t?�[P�n3��f�w�#��C�P�8��Q�T%2�i��U�|�F����0����`ch5�e]����@��+����xJ�9�|컎�")`����ճyd;�-t���Y���>n��p�W'x���_���w���ʢ�*�q�P����.��A�Ƃ��|�i��ġ�͵�����T�{�_�k_�sE��"��i5�7�����(�*K��IֵmL<��͢�/��FءV�T�%?�2�D,�%+w�y�c{��[Vտ+�+/N�~/�p){�'�:�����LY�+k��k�J>�>�����H����ʍ_F���=�q[|)�G�Կ����"��L�n\�R������Z����6�����$ߡ�ש���B�3s��J:c����~zt?�g$dkaS�[/�[�}�Kq�>�q\��࿘<��U��R����_�ʐr̍Vs~1�&���ㄦk�D� �6�&t|~�Yt�E �������=���(D�A-~�73��_C���r?�<ŖB�С��g�*ǜKǹI�-@Q�D�ڈ���)��i?��T̀��<*'�fS�@��|~�jo�UD��e�9ڍy����%2��KC��R�W�@�4c�[1���!�*�`DSX���V���������J�ogv�F(S��i��$I��Y��c��Q䓷����D�e��f�/O��#F�q�-���Y- T�P���ˊ$\����R���!�����;�-���M�·a?I��^�|a�lR��yL��p
��&nl����i.,��g�k�N��#���MG���d�n0w�Ͳ7Z�G��I���\�B6��6�{ӹ§~�s�߼����7u�
����1*?�ȷ�e�`/�<�f���~��D�1S�a`]�Z]p%YB�F��GP�L���ۑpo���i�rm׾J���/�!�p��� �yi�	`NF������ej$x�L��tC߇�vN�V_��9��~V>�Vt�	�S梯�%����Ű����^�E<���Zv����EU����$����w��sʂ}��7�Qx�r �b8�Vκ�s�Ȩ���e��7VrN�8e%n�����'���P�1��ϩ=�@|d�z�x�o�G��.��� �}$�I(@�1�@�����/�\�Éb��$�l���V���U�3{���JaU��W���>�	�d{u�Ԓ>%C��m���r/��&�O�����"�	e\'َT	�����/6
�W�}�[�����e�g��0��J����מq���> ��2�Bʍ�
�$^1��W�UX�d+�4�v4�7��])�=��n����$/�o֞�v�?Vº[�
V_�T�ˬ�4jp����]�eRZ�-�cR���k�B��ja�5�����@v�]H-ηza�r2:G��\��yK��i0���޸$J�GN9��e��G>�r,B�o��9����3��9�T��FHpr��Z��C�1�-�~c�:H#;kFQ�]{�gSC�J.�l�A\5�Į�4�w�{%JBv~���u�N�ePyk�<��9.�i7���Y�ȀH�]�+-��K��;��Q�k7�6A�N�������h4�.
Kl��O�[Ǘ�8��#�.���W����=ݫ�ɂ����-:!�0��ɒ�ja\���c�T�&����2��@�>$�Tg����V��V����n������p�\����qA�bs0R��I�|�*�0٥p��E����Fa�^0�zE�}�ֹT��[Ȩ����Hw�=2�$��d��� V�">���5v���P���� ��c���FF`M'��@�[z� 2^�D/#�����F|���7[,��?lP�z��J��\W/����FK�S��Y���44~y���-���P��',A�.����h	�A�������1J���1�����i|`��V�����H=��A���/ki����_T�*�c ���}7�.w��[���E��]� �.�d$�O�{K]h��h8�����==��(����� �����,SH�|��`��n�ͨ����!A�O+^�OyE6�3��Z�*ë�}5���D|-!�*�t̸{�B����n�����Mi<#/jܴn��ot�)�8��G�gFms3	j�]���&�iR����S����/�"D�O��h�
����(LW4z��FF[p��B�ߖC�l����۲�.V��gvH���2j~g�eQ4N;����%ْ�+��+˜p���0[^ow�uNݝ��앳%4�߼!U���h�V�����/�ٔ��/P�D.aq< +��(}Z p<��y��~3�����F��C��i^�2E�k@i��%A���Ōu,Y�\l�啊�B�  �w�O�2k�`%O�U�6����?��_�Q�s�)0y�C.�&��z�@�M������N�P�h�TF.	L�HK�ŻDf�vi���������*��<���W�#��8F��M����P�D}g ���6!�.�!j��{ｋ�D�V���k�轷��GYK����X�+����_v�9�̜k�k�7t�2<R�wQ8�왠��V���d֛���}R�y������dϧ��%����k5��22X��~Zx���,�ubN�)5�Iه�}@Ey�-����L�Z��R��^���ȷ�w�q9���;���k%���iS8�����h��4�͊��*��yW8ty\>�C�9qsN#(�4U%����%O�-�C4	[9�>VʍG^w���B���-�(
��ͣI�xu�R^��(w}Z��И��B���2�%�"�<ӵ�$������Epn�k��(��b�
pm��1)-��U��nk����w�	Z�c��9���ܒgA�2�����ea�� o������RD�5�0w�a�J���(1C�e�/���'�ѝ9"���%����p�\�y��/k��s�w|��F:��4hǓ�'rq'���c���7'PF,[�Cګ,�\����=o<��\Б�?͠��I 4Usu!�W7����^��(CMqľ�0.���Q�[������O<%Gr�px]�����<�P5��L.��!�[��I_>*5�O�}!�u}�BV����]?����n�w)c|~���Y'IˬO+)��0O~����/�O<�8�a'{S�T�7�~��덩�W�m%� ���Я"
����t�	���<����E��� �6��s�n�&o󿀼Ws��fd���l�u�{a�+{窾��{BG6#�R!s��.д ./���~��N4��!D8z>뗔	+�E��Ԇ��(r�"^��7/jK+J���|*���@�Y�O��g�m����yH���h�4˚Iؤ^���F���Tt����,�*������"^A���"��?�QkGAb�Gn�������FB��MC�H����]��s�U%y%��Um��W�
>���O���'�6{�,8k2}����@�<��S�P9���L������eB��F��K��	P孈�Mg����za^藶���C��2�A��Y?���U�Zoc��8��:8# =��^ �/��g�2b���������Ž`�阴Ư���_���[69�(7�r��˪���Y��$�����;:s��6�wI�|<ُX�7gF���?�|�k΂��JU	���U�[�8w�/C�K�C+\�����ט���Ž_g��4}��BKg>�5T-|Q��7���Ȳ� ��M���>��Eow�('����#�>r�����R�~����� ƺro|�U�_�'�'�drƆ���yg�$Aav���U����3\_�g�;���o���LsB���[-�l_�F��ZD��	�ϣ�v�T��^�Z��ȼz��]��|Y�2O0�aYe+��v��E}���'ѻt�V%�g��A/��1)����
��~���ݐ҇�w�~��Rk(��+��ZR�T�ǣ��κ��_6^�I����i\��Mb����Z��G�����豧8L~�4_�~P��uV�K����nw����L󭵘��s�<uf{�����]�� X����Э��a�iF��Ҵ��-�[6���V�>9Ր�|��`'��)�Z��	�����}V��,����a�5)���Z׋"���W�\��)�=,��.�gO�!@�����i�fTMr�v+9��{(���5��!���Mf�@�)⨦R-î�,r7�%��$��:��B��J�x�pnE#�F��F���m? �n
���X�/J��� 3R�Ͻ/�v�͐2�Q'e�Jʆ|�O�Pc��
�ł��Cˇ�=�V�T�
����	�?����LW��/OF�0�y�xOTe���a�
����`�U\c���ؓ������<���v�J��pe6����mÔ�V���Z����e1ԉ��Mzp7��Q��t�'e{��_��Z�^��Ӊ{�Ŀ�À�K��p��HuQ�@�� zC��*�Bye}��B�;�I�k*K���e�W���k�M����=��
��G��6:a�5J~J��G"�W���B��{�F�fi����L@��~׺���$(��*��T�O�״��n�u��O��	��%�ߚ�W�|W{M��o�OhS���+��}���/6�<M�⾪2����!�v{�qnRn_�t �����X��:}���#��j��� 8�*/�mSN�2Mޕ��g��4���b��p���|���7��h��N(Y-���f~c�����������#�K���n},w�5�t/R��8��y��k�+l87�ﰸ�G�!.��Hj�ν=�����1S��0��ګY��0L�K�c��E����?v6��Vƺ!tY_��D3��w���$��*nL��i�P �RE��j�}.��E�i���ެ�����nf��RE��W�=L��UUy{N>� |*m��%��)z�΁,�������v�F��طU�h�8��$#Ջ�~��t��l��:���=�9�� �k�F��0�2ǒ+�a�ν۫����y�����/x 4j!J���0:��ذ�Q�!��r��'���Lӱl�k� |k�v�2���XO��|'6S�+=�̒�v˪�n�"О�~?O#- ~�_k��*Dx�@l�زb(Si(��*�O�(Gp�c��ɯ����HP��oW� �r=e _�w�@$G�(����"�;�d�T���ӻ��6	up9S{���4�]_E,쉊���l�`�)+�!�5�pF�}9:#ⴜ*eE���~P��a���jZ�����d�������̿7]��W�i�7xG�TY�5�� D����5���$�Ф(�5�^R�g�J���j�&.OQ�m�En�𙅏������F�$�/R��/�3	U�Z��'p�FL�g�z�r;���mN���ۈ�('�f��%�ڡ��Vk϶b�S��4d�)����H��=6��i��p�ȧ�.��.p�'�b����C)��Ȧ��
 �O
����0/ձ�bU��PD�i�3E��~���%K�NC|�#�YnxF���L;��`�O�ګ���Rg?�m��wTk�j(�WE�fL6��ؿ�(v��9��kDː&D����&�߱}�h��N�\��/��OX`S�"#xu��&�QN�Od�W���_ <�].i����S��Q_G���0=��>�Dlo�<�Đ2T����~�){��R
�4l#�M�_�ZPT��O��8�A�jZ���:�V��r�5X80��QK��3�Hd�����A)��?�Z=r�u��ܐ�>sO�zqO{��:�ǽUq��w��U��X����Fgk�[��i~��c/q4�iF���m5�@0�$8/ܘ�n(c~s���;�c�6×��;������$�-�P'���CA��b����_�������_�,���RƗnIs1�κ�� /JӖ=��)�Ď]��gV5�q�@�%qj���u�� ��1h�-�X�j3)��W$
Տ�@ �Y*Xӗ5Pj�Z-m����+W�{Ru��l*�շuVX���8>��ϧ��&��o���w�������v/D62=��\;ę0��<)nCN?�a�洔��� ���7콩�t�	�d	����f�%,���m��Y��n��A���t�E�ߥu>��-�K��Hw�a�)Q���*�/O�������o}�W���s�gқ,�u[B�M�l�0��d���t`�E�����ߣ��g��o_��Z{����~�Z5�l�0�%��S���oØ��$J#�=Օ��D�_/D�zD0�R�NS�#X�,��ƪm�^�?��(��0	�����gy-�����|oK�!J_ $gJ.,��~]F�0�Y�"�?����8�E����Q'COz}_���L��V���{����	5ͭ6�-*y�!��U�a�N�4�P���	׵��QZo�RM��*�d�� A�V$>�8-��//`�����2,�� Ѫ��Vn�D��cK����U�k�y��q�̝x�����)σIӡgʊ��	A����(z�F������^�������#=�}��j�H�L���P�0���=>>�t�Fӻ���#
��	&tD�|b.�2"
���6i�����pVV�q�X{Y�~�y W}�[*�[.��{���Y�f��F8�m�M �Qp$aKo�ݧ�����{�ݦ�h�\�#�_]����ʙ��Ͻ s;]v �<���.���3��r��|)@/r����`quG}X�{�_JЖy�8ED��P�kE�XGjk�L�i9��AN�ǿ{$:�U;ś�#�wDLQ;[��I����K4$D��^��r�u4ҽ)%��|�����g�OL��0Q�=�L0J���n �yh�Ѻ5�ɌH�C��dt�6�m8�Y�tTT&����BU��İw�&�^��9O�-X�UD��$�\��PK�N�f U�R�o��\e'㟻\��Z�{��E4�4R
`):4�!k�^}�[E=�S;�(��+���I���u�#�(�~�@��0��<���7nFA�&>.��#i�GAĵ���l��K�Ŗ�b���T���3�G=]W������X�ʉ$,��ړ?|N��}�m#��&��5۟�#�;�m (�7�US�<�M�4o0G�����t�B��rvWL ?Մb�Z�RH�s��x�w�z�x��MA���*m���|��]����G�A�/. af��ʇk��ͯ�z��E���a}5�^KԚv���{��~��ֈ���bp���G1[��܃�L��5�+ϼfJMe��d���T�er��3����u��5�m�雽�F�h0�b7�P��G$m�q�tfyI�����uP�\�=lr���tX��ɪ�H[�
�h(���r��b��#x}�(�8�6���}DG�G��N�`���"/��ֶ���!ZIx�߀�3m7�!�.�K�GW껊���q��z63�XW��ס/@A��A/ۭ�/sNn|�Td�l��[#<ެv��������,��a�7k5�Q�v��3|ū�ilp+�S������T��)�v|�2]��
-n��C�s��F��:�)�@yʊ����C�4$lF|��������iO>F����a�ے�����+8�3��� ?�s��&vm�X�S�W�c�ʇt���ϲgn�`��d�?,�o���ƾڟ��j3>K�%zs�`�{���ū������1o��s^�f��y�Q�7���rv �ܲ��G��`�":�Ĥ��[���-���u��������oɋO#D�@K��8��^��w��r8d��?)���y�^���ܱ�	��,��_	�ϗ��H�S|��H�k�j�B��K�v=�^�33��u���n~n��4�����s=/Rw�ɂ����}{�fvE���#Y�Fo*5Z��gr��n^a�y�����v��сQ3�m"�p�_���Rq�: Eym�\�p�J�qE��Nm����L�޸@.���N}s��roM&�;vk-.�B�D���gR��mi+����Q�6�ﰛ��1�y[���xg�AFF�TNs��!N�$"A)��&?��E"2����M{M��>?XC������M��Zq|���"�]�;ov��}_�o�	so�o��=��O��T��.uR<��p¥��:/�#��n�}aT^ضt�^�� ��R�k��๗Y%&x���m�#��ˣ��s{��ܑ�6u�q7oj�0�CD�L�|�umi�������2o|�^W(�>��+���X� �z����s]��cO�c�F����]S^�5����5"R�X�h����-_��A�jA�:��7x���q��ջ	eUr��0)�O�er7�AN�-WBOy�ވ+�"�ߥ��dK��� �6��=�y���a���}�qՊ�{��t���~��0Ӛ�t*��j�CQ߉8=�Ɉ��g��	TQ������o�-p���1$\b�߳��ș)���h���C��~�՚��;Y�T{	�o�,Y,�[=Ǜ��D������9� ��ǥT�l��œPoڮ75�i��T[Bz�	�����GQǱ�H ��:a�`�eȑm�e�qd
z&~�=_����Bx<^�27�m��>t�O�g���4%.�B�r��#��{o�.���{��#��Wkv�RȌ}�MHr��ۦ?_�cƳ�X`�I�����yB�����{��?�W��/�	���}��|w��g����v�L}�>"p���ǳ��qh{�g����»]`�G��Ae�:xW���iiA�E�)���{�L�k&���!|Ķ�)���,��*Ο�|�n�N.�@��+x�)� �&B���7v�1
ͼq�Q%&���[�� ��� y�g��|�<�򗀍��l>�Ҥߚ̻�q�]u76ߡ
]A�ӹ�?�	���$]�ۮ�fi����4�w�t���6<0�q0�
�B�����=��ٸ��U���d�egk���
w�7��+��ո��n�I����x��J��榞����i39�}�lk��ȶ�ĭx�(n�e89���»�ns�͹���#���K��� S���]�� Y�nf�8�f�c���W�[ e��;g�C7�����A3����;�/�Ã�4��������߿�~��;��2'��@��K���H�t4@w7�0h/G�yS�hZiZ�����I�K���n��=�7e����:��6�4;�́M���~P����"I������8S��EViu2�(��F����B@1j��j-.�� �M'Lo������%>f��1&�������}��1}�/�=d�|��o���C����� Hi�p5���j���ڥ<+q�;i�����?�U��[0��W7�Ov�9O��A;��jE��@c�<�Ҙ-y�>ֵ������wZ*'�ޑ/���}���[-XD��Jy�Q���x<3�
Y��`Ŵ������m��0�f!�]��	u�t�cYA'�M�C���Ϳ8c`�?�=�x��r�;��1���ZI��$�p���`�u�����ؠ���E�GV(�	�wu\�a�����#� \�Y8�al_:�����&�ݭ���}�}�Wۭ�f�i)�oaÞ@_�Vhn�;���b@�Ṅ�a�E�V��x��m>���H>�Pj"���D�so��Mp�)+��:IOdh��a���4��#c�pl�o֬�x�]T���$a�$.c2E_k��G������* }ѡc����A���������K�V���l°�f���Vg�q]Y�����琔���afu��`���O�%�5�ټR������8�����O[�ǥ�9������*$8b��2��I�b������3ݤ'S�^���u���U[�^y9ܤ�v�]L#%��"Ɠ�t�]ֱ{�$�C̽P5j�S�����r����_��,F	!~�&V�=���xj���c��c)�50� �ğ�C�F����f��L\jA���8e'@,���9He��S�`d��n8I���P|Xʔb8}��*p?���stX���J=�;�\1�]��L����h�A��j?�!�����ӭ��Y�m�fzU���3{�b�H������~K�fƑr��T��	0�,T���bH��C��K�� ,���A��ٝ���ŷ��e��p 87A�� ���TN�9Wyʿv�I�K�<zE�ȴ���X�:Ͱ�p�X�C��~�Ht����}�nv��a�SM�NPN4V��BG �J#=��T��$�0�箊Q&�vgĚ�}�G�����K&p�4�=��@!K0���C!�%휤��>!�ڒ����Ѿ�p�GT�,�ae6}޽ot�3O��Ŏ����M�lG8���4������3�yV� g�
�� �X���I��d�����Y+f�!Ì�|����ӡ?��j��U�(C���i�78�{���+���I�q��S���UAX!�G�P��6�\��_J�)��_���s)���y���x����u&�CV\̫��ɟ�L����1�#
��*V�o\���\7/�r읆!���Q3�-��q�����1�8$���y)�i1#��}n���Ni��<1��446�/���%E1��8��Zd>�H�qd�W��ǩ?5�8%rOv;�����}`��nʈ�Y[C'o��Z�E�
���li�x�,�d�C���i@����dO�HiV��J��Ï��zǾ�Y痥5�s��\]���H�'�>ƌaB��/M�q�����n� ��`�l���a�<��`������!<�	���i�������:x0w�D߽袁�O�Z�WpVE[�����^�3�X{Ɲl�z��R�^n��XV�s������a?�+��Muw�.��_�ˀ+��'3N�ɪ}��@�N|�/:���<�
7
꧶�OI�2�����7��h	�?d	_V��g�J��2H�>9\��^�&��\'���̬Fy��u�^�׼2��Mt���!7�0D�N�i�o�O�Ł��jIR(�@\u�	qg��kb<Ϫ��봎�7���m�XB�m|����Ƅ��s<0���� ���%��?8�������d���)��Q����s��aǵ���029��ӏ��NV���� �grjI=�˱ �ڦZ`A�Ǘ�8��zLM+b�w�4.kV�d�Ϥ�n��&VŢ��ghP��w��F`]�/j�v��o�V�I����Ao�/�|r�{@��B���a�g�`�~p&���Ԕ�'6Њ[SvƼH��P�b�|�*Nk"Jb��˕�i?�ɋ�����ذ7brK�j��Kׅ�=Z���K��̓Gw��'�W������jA��	��i�B�t�d֏b5�OMPk��]�BDp�69�*����V�U��q�Ŷ]�>�k��ėg�*�HΗ*\ W]6��|�/�'~Ђ7�9Zϕ9P�W�D�2O�5Xr%HgΒ��i����_�u5gά�f��i��*(��8���K�9� �X{]��!�ՠ�����[
�ʷy"٪>��TV������҆��lEw:��:����jr���tu'�:��qMa��=w��kg��k �t�X�p��GN�p�땷 ���a�9��M�;�w �׷#�vu&�K�
w�'ެg��e���1T�<��3��gt�4>�l.�Y_�7{�Ij,�P�@HE��NxOl̰'%��4|^�P���J	�B�f%��H̳B08��t��"ri��#{4�/�}�\d�(��d���{���j��O�8�,�i�n\ �������=���h��/�΋�P�m�p�6�&�R�O�x�Ja_�u|�ڠ:<���F�R�@�?^�ܭ`��n�]���
8�)>���`%t:~2۴��,z�lg��(̿�#Y�������b���v�.�w�����R�����Qߜ�R���t�(�@��I���]Dߺ���=О~��rG�8HU����e�i}��-�Q��8��P�%�5�(��� ��j��+�O�I<�,�,���50�z[�[x�$��z�JC�*�ɒ�mP�-A�+��d��{�3*dL�0�_v��-���z��T5�z�����uTq�.��K���}B{�O��.���G�r2�(MUz�������|0�G߬��QL�{W���&��ťBi�l�߹����Q���ҧ�M�7������=ت����tT��p��] �M���_i�����wH¹m�Y��%��"{�I����F��9��4E�>'C��BVC�T%���O6����]3���ﱷ{����y	��(cW�F�W��e�U{�'���G���}r�����;�[�/�o{wOýYC���Ga%;]G�M�C�Ǯ�?��)���� '�3�����F��{��!��Z^)6��=5-���:'�T::��D�.ɷ�3h�G� }�K[hݷK�#Ϳ_�V��A!��u����&]��R03�!?�:����%-'@�K�̾a�;��z�����F^\��&�Yj�_j��4���h]���Ә)�^����iYwvO�L�<n��~VV��ry�����^,E�!;��W����N�46��]��v��C��EO@�Ot�t����N�u��L�ب���ߓ��2�.�
���/��<�9��E;J�b����"�e����%�Vo��9S�n��#)�B�CG[�G�ד��]��n^]��7����<�h�/ҝ���&Ý
n�gS�p�x�߳췏'�ճ�=�q�aV�pEV���[��ǆUbt*ag��R���0������/+�J�h
:�6�s�<|�e�-�Z���Y��;&�;qL�����r�_<ω`�R�E�Zw���t����N�G��'�E�&��+�c��Bs��K�H��Z>
�`�o��=�Vi�٨>p��n*���_a���Ҷ��L��~������i�җ�n$e��J.����mk���W���ȴo����\��GA�oҧ�Կ��x��0
l7׃�������®�� \D��VX 
-�+��=H�8E�$D�?»��5�6��uq�Njk�
�W��S/(%A m��O�uJ%�±��:ծ_R!���@�#�><I$��5�8]��t�s���d�#�<�屮"��U��z�+������.p�^I�q}w��� p�cj�Jp^�K�P�D[���ă��J�V��-	ؐ9j�˲J�'�1������Mg7$�Reky/ZUj��Sx��D��Կ�)��f��0W����ʼ\��Ț9w&ѵ�
_�������6`	�����*�u丨	QX!�nɼ�,(�h�*B0�#�������z:�k �hȚt��\������m��xn'�j������ܒi�L��g���l�7���4gWO$��}�||p�;H?-��v��M��� ���_b*,o��?�v"��x{:���[5��V�;.'t4��,�)�*�������7yպY��}>tqS���H��ND�9�n���ۑ�UȽnyg7�ԁ蓴r{3�/�`o������T�W=��oůF�)��7i/D�8n�ڱ�����l�n���&���
���N;t|����+��T�Z�b#���G
m[���{c�_]'��\6�����6�V&	���ͧD�7O���Z�]�u�7Kd��Z%e�����}a�Ԗ�Qf��T������~���<���'�)?�^�b�͹/�!*Kf��w6���DAp�����zh�5Y���B�w�~K�Om���!���G�xh�8{@a6�$�T��Sl�&�Ў�'a��ထ��F�7}Fl�d+j�܆&�mZm<НC��E���Y	5��d/��������[A�f�x������i��>^����p�~"��\��N��������@զ��
��lD�*�.�	>|�7<L$=Nirii���m�� ����v������ͥ��o�)E��I8I'n��Hr�v&�:�ɒ#�+���#�w��6P��|bd��Jc6Q��}�ҿV@+�-�26���B�Wg]?�y�-7��\�	*���tqጹ9����Mi�{`�x"����d���$�-h��X�sw�
J��F���l�}q��Ѥ���ї����Ů�]�:G���M#S���yg��_&$�+QWZ��&νjZ��H�~N��5�HX�a��8_S8����X,��X�9��d˥�C��"w��\�Pw��3�́��lC�����@�!GW��m&绊�w W�Yw��[���Q��*;��(��p�$@���_�
Ӟ��59��GEᤴ�+��8�����%�����;]�����On�����c�Ϟ��/�]��|t�_K7M�?Y��g�9�/홭�`�;�W�W�P��yԚ؇�7%\�w�'��}�4��x�����Ԓz%M~�AP9��0tnP%ȡ��j=�4�i����)��x 2��h���P����N7HJ0=�N�ZoÍ����tnsq )�"2eH:��
�x�Yp	�0�����o�t�VRdh��;V3r��ry�􃿶�E�]���΀sR]�&�K�#B�d�j2������?�`�z �aX0��3<\͓��`Nʥɵ!]<W��;�|OPL4� ����s�W�B���~2j|rvX�K*��Rk����.c/�3NQ&)y�.���R�	{7G��e���+��"��%��=lPJ~/�@�->�O�W:o�ˠ��z_G3�'7p?����ó�,��ܚ����3��IRh�F�Ћ=p�"��m����[x�"h7�50&OEL�#A{��0���r9���Ѧ���W�� ����$K�F^���ܣ�(�hĮ@fiY���8M����r���=`6��#O��Yd�5�#tܝ3tQٵ Q����'�@䳇���������`���L��0�wN�I��jk���2fVA�,V=��}?�N���A�;�K����`T���=YYB�шro/0e���0%�8�7f"�^2��u��h�qS~�ji�]����w͂���/α茶Z��| ~�����Q�:V+��g,N�.Va���R�pǿ(.�x�2��G+��Q�zi�e�n�NO��'T�=�&7�{�!�nL(��f�I���%�Lo-��\Ҍ�6گ�t��W�ָ8��R�8=���f\���Q�1���h�-��-(H;\�G�:]���ٱ���;�#Q1OK���M,e]X"(|��=Ĥ���,�����1�_Y�I\��������R\�tl�f�t�r��G�����Q���$u1�l ��y4"�q/�M�"�h��>K����~�Y��/�n�(d}�iΰ�bbL
S/R��l�.R��Q����N�l��(5��F��wßcS4�5��/���_R���9��,�R|A�|LK�Ǉ�f��g�����=�'n�I'*�M����.]L��Vȩ��$;����
{X
"��*����VǪO�>�I��U�)L�����d����|���g��G_t�?O`�i�����vPO/�c�]�9peO��8��?7�����!X6m@��]"k�<?�c��qˢ����H<�s	C���w�YeW+5?{��D;����2����4�XI2Q�oL�'Ih��
F�m���l���_����3Pe���b��*I����E��yaF5Q	4��O`P����7lu!fݦb# ���%�ɑJ��
���z�����QE� �I]&T�r��I
w��m׎\y�q�w��;]Ƕ�^��<:A9����ܤ&�&4���{]ဖ���jǷ�Ԕ��O�S�aK�����Օcb�{}U֋���0�N���p ���03O��֊"�,�:Z�K���tӁ,�CCϴ��4w��z�/��l�Y�@w쮝�z�(0U� ���h��`o�Hر���V�뽷���Gd��x��I��^�H�ڦ$��|?�{+9V���m�Дh����e�s��Oe�r�]�I�7%.��<44�B�Г؉��Uٕ�.Q�����ͱ�HnD�Fy�����x4���Ҍ
�2!���ҥ4��֭�ї�H�R�����m�7��{��X5,�O�#s��n� z��2>+��i�80�	��ֽ�Mu\	�mW��^n젢DG��~Iq� )�q�VY:����9��rOb�j��}G�ǐ��_hᕸ��L��sC�wy���RW����B
���XKvh�+�"q�#_��C��梟�TUX�#9��Yr�s�?5D@�:�^iV�E��qh~ŧ�nت#SǃV+�)ޫ&(A�R�<0�2*wu,������I�4���T��^��t*��ȸ�3�I��Z�H$\�Pf�?��X��\�,P��ց�y1��;�Q���K����.;�F�;#�*V�@_�p�H'h2�%���T��,�l���x6��2�]N����m"cD�/����>�낌j~�6�Q�Lw������h���T%�q�h�u�	1т�
���.$���ˀ�fp�ki��NѝP,����1�Ϋw��uON�S��wت|'^M$����i���DӸ�E<�K�1���������*MN.=�_��d�A.��I������ϥ���{՟��;��J�\z�� ����B�|��~/�gG	�G�}0�ǖ�����sLW�� �{��5��GRDO7�9V��l9z�> ��6�~uw����l��������ZXa�h�ޤ�`ٰU�o���D��������݊.fR�;�[X#\�lZ?������^P��U�K���kq2]���������r���Qұ�K�^���OD}����X3��L8|���ΰ8�m�;�5x����ogN�]��H�$T�M�y��E��O}�A:�"?���|x�ǖ�P�G1�~8�[, V�쑰9<�F6�؎�O�ϯ]WW�B
�!�\?�t�nĹ_=^�}4�^c��G����ۇ�����_�6��s?��wv_�m�B�	(��~ڭ(D_�����Y�}U;�.���胦cn �s�a�Օ��p�V���Z>�,�^2E z����N<j:�����P��o��'⻺�q��`�8�T=�-�;.?�V��$Vs��ҼG*}���И��N�Q�Y��e�\�49�������x�;�[����{�\y|֢�j�M�������U'�V�F�a�Nl)]�_��H*�^+T�%�]�=(�s��d}��o�s�SW���f"��(��Tz��+ ���O��J�>咀��Πp�M^:�T?Aju�rǽZ��bݻ��c��]�ԈGQ|�<P�����cݠ0c���bZW}��j�7���=��Yt¬�Q���֍����3�v8��ۗ��G��w-l�������eqxM$N�p���� ⽼G\؞�l�u F��ri�K-���O��5��-h~6��
�Zx�eJ���*������y�w�'0V��◗����"P�t�Z��<�\��u%�D���Bp��NoM���q� ����k0�c���
F�T�s���/�[���Z.���1�k�M'�a9���>�[�S��륣/�V�y�U� �s��7�x�/a(��#�}�e\�kdJe��;lm��8��.�q��fu�5�H�Sf�,r�;13IJ9d�/�j4x�9)F�k���tMKܦ��s�X&���7��ɯ��)�pS_�F���Mz(��0���/�5ݟ�A�Y`��"�[s��m��Bw}��$�A�S�ޏ�%��3#oi{[*\�}�,��:��|=�;�����~$�+=�pڠ��������~[���˥��D`�� 8��{��V>5'Z�y�76���%E����8�$����
�'\*���f���3F�ӹ)�#x��ceq�y�]>�7Sj����Vzy���=�A���yZ��"3����LER�����'�9vh�Tg�s�|U_�������[<��#ȑc�6��U���r�<�n	�"�B���6�
�ç�����|T����wHH*%��C���$��1M4�pO���p}S�~͆r�ŷ��;t���
	��;��<Q��
̙��'���FzV�/u*������q�/�մ~X�(��^Q͡��^H�`�hMzu�3L->�/���KD�����v5��-��
��^�DOelԢ��+U�~y��s�0���n�� A>�j����|4�<���X0�vG`z ṲJ�`��Ð��Jb/�g�@��ͻ�ߓ��f�4�9��������+3&I<���^�){G%�0P��vEٍ��ۀ�o��:�0���K�i)��F��
��U�LI���ՅNL�,㰙�J�cSȮUe<�a��8&�5~�I�9�y���{̑_?�Ъc�V����k�قi���<����
�GH���z���s�H�®��؍[|�┧}�>,��r��P�hFђJ�'t_z}����	9OӉzrA����K��1E�g�I�
J:��'��R ��z����~p��%��C)�-ӻ}��߹��?t-��ތ��)q�H���>ȭC����4�R��1s�c�r��B�6\��{���@$ɣ�����.@z:����)f�o��g�W��43���Z����YJ�oG�ئ"v|�?}�th9��h��/��OV����z_���O�E}o�J�t۬���������[A /�>��p���sU�{A�r��`�h��$ۮNj��I��ZEwr�&��vwk`F��[4�-l��s�J�����s���y�N��	v������I_C��xV�ՙ�0�D�����O�ER7k$y�V���3��
�y�Ϝ��՞
6F����^�z�wF�5��ⓘ	T�y�}��7�m^M
��ʩ�۵��`�p!$�<(9�;;��A�$�l��'��'�ߘb��+})���º�����`9�<5�6�����8;N�gP娻�V��E��vmܘ06�A�H�i�#F�C4s����Ōe��ƨ�zG�h&'XN���*�9�a9�.X7z
�;BD^���_�/y�8-܈v0lC�"G�g��,0
7����SM�k�\���V����V�������������B�rq`�妱��I���(n��p'��u�����!T�O�8@��L�D�p��k�J(�]&�/�|����C���I��'��a����nF,*��/�n�x��;w��ђ����8��j���e��<��OJ��}�ٶ.���ʨxY�����M6�^ ńtX���|������, O�/��bLz](�VԓĨn���eON�:�R^]�h=<�e�[���R��t���M�W-xE\��]�a���`�Xːn��&��L
���_UC͏��j�������oQ}o�(Hw�t
H7Cw	����tw# %" 9�HIw��CHHHC�H3�٣�����7�k��a�g=y�k=k�p����`�X��V�b�}⧭� �P������lƷ��I:#*�SZD���Z��)Z�`���.��b8����k���A�͑����ѷ_�op�ō��ln�u�"��0�\*��9��Λ�>�m6c�ë �'���o�Fƨ��=i�wÎ��]�|�s<�4��Q��\�O1E�i*�����`Z7���CA���f-����D{�L���ĥ�)���~ێ��-ߚ�WП������<f��onO�L�OZ����"ʜ��d�گ뭂��'Q�n�B;�*���!��A�'m㺔*�z-]���
�)��tx�u��8��1����m1B��b���#�>׉�����Z�p�=%f�P[��"��YH��fh�^l���+Yx��92���e��U:9^�q)ِo�NJ������I��Քh�Y	�0_�?ɉ�f����a+��˔���b�z+o2-CG���+���&l8.�`�'*�E���x9W�yA���j�7^ES��F]	�K�cu*L^0�A��¨�B2�Ϥue��{�VB%Tb:=l�p=do��j_���]wv��j�H^��G�`����P�qx�<��˦܏S�2�ђ���O酨��[�!5\������U��<�7�F�*�R��N��M�3f����5��P4v������7�����DiL�8�O�W"^�v�7�䆋�� ������Uo��|#�~>�G�FnL�����A�f���������@
���S�-U�X��ͷ�w�G�Fn�w
�Q!$s���.������ɼ�5L��d��l�+��G����P�얫@�-�ܰt��!c�J�����"���1C3��՘<Ön����K~���L:@-�s�6�Ow6�f�o��F�yv�I�� �C�׀<[�!>p֭�����\y|r>��jt��r�K5��:/G�+F�B���}�W�PO�-�ũwSE�cl�`��΋���GVA�3��W�S�Z���@���5�ikl �W�Q����nV��쿖p�x����j�����ͤ�{� ��q�꿨�l��,����U�i��5q2Y����E���%��+{��j�M�#�pJ׸C������,K�'
��~�)�>O��"v�ڕ��%��1$^LV��lى<�X��.�:��>��iu3vc�g�W6ȭE;�D3�i��VE���>�7���K/�	ӻ;�3�/ԏ���X=u�¬�ꃟ(���Q\��d��q��z�U�-<�J�P�->�tOK���5e�D��\�!�� ^�$���*��3�kUc�]�3�S����͢��r���-VV_�_f�Z�d6k��@�q[K������SkH��?О�'���D�3�{��������M��&#2F��"2�_��֋��i1��_�
H���r���H-�qj{|���ԴEA�1o�F��Ǐi�Tz$��`^��K�x>����8J�~Ɠe<���`���m�LC�;�@�_U�l����Xo��>��ۂ$�4��}��-V`s��v{w�ߑ̄�j-� ��jHz�k��q�.�HC� chd�w0�R�~���o7�Z��96�i�i9u��V�N�C��8�N��v������&��|��;���R5�[�^���á�����q��U�q/Z�$�><m}���� 2[��_8���i��3�?�Au���� ����I����jB�z,[rg������Ϡvv��rJ��jS�qۿ	��`�@���f��cXx���g1��Ѱ����;���T�Е$^��d�,_�K��}�s�b[Cq�G�t�.�f�wt��tF`�`�Z�� �����N/]D�.�U/�=D�(_��1����(���8Y�;���g�{L
��>1�?�6�Q�1֘��AM6�D�v��e4,��7�, ug�g��~�E�ZT�p �%n!��j��|_M̮=����D������9���`�翂lI��{�L�"gɒ��4O�cOd/�Z�l���_8VfV^ַ�od^�ōq��#��f̈́4ʔ���lMX?sߞ��%�yӿ0�؏��9��(T����H���c�� _,U ���K[�ߛ`�783p؉�J!!{-,eo��G�g�J��]���3no�B�Gݭ4)b�0�Y�6T��^5���P����)�y�4)<yO���q���C�m��b:�NO�;����g���  1�$F6�?�zRz N�z�!ہZ� �����|*V(�������� �"�3B��n���o�`(��9��U�y���@���U�ZDz�d��Z&�n7U��������eK��B�wP�'>�{�k.���E�.�>.���/�s��pk����+P Nt�K�f��YFr���q�%��[��<��@e�E�X-��?�s4���	������-~�>��ү�'y/?��1��3�� �N A���ɂ w[��>�C�Mƈ��u�����Hw~uz��L�J^~R�X'V�d����K����-�8��Eѕl1/�A�b��#ݪ��N"�҇B[TO~nR�1���CJ�~6�����8G�ϛ|r����.���b�����'/����["��{M2Q���#J�p�U��2,x!��h���Sř>?4�eH��z���|����6 �*���)����:�m��Z�Ь�������D�N ^	Y�%~�*��k����8'�g�d�J��O�XSKRv$*Lmo�Yt�ʟ�|X���"�v���eT8�����I��&|(�l	T�A���t�r�x�-�=����ώ��)3;�w����8��ǥU�I���-��
�I��8Ǆ'S~���3�<���N�������Gc���ƧR�,���B����wL��dYg���xy��jI���U'?T���.�Z�o���s,��f^c��،r���˚���ȕ�nI�;/�R28����Z�1��W���^.�d��M�mrp>~8F!왕������d�n;�D'�p��iZ��������t[���\�\?L��	����r~��V����x�������������ר�X���}ɩ�F־�	
!�B�lR����Zp��`[��` �Dϕ���ۯ�y=j"�b�q':��7,[��Vab����1l�^��@�j�{6�[�s%վ��p��H�⑱�����=h��"q��@_�s�0'�	kw��O��j�0���A+h�5��3���>�i��C�T�Ot��k6�Ζ��f��Ȉ5��Ơ���ZyA�ޚ�aY�e�a'D�r�")>���$�ZY
/]�o��Y�Fpm�����1����O4Op�=O2##�*�_uh=p����'�g�;���L�\�N�)t�u�c�+Ӛ�8�+��ఊ�]�h+�����9d	i�� g���( @1�Q����Eט e�I��Phoҭ$����[u��>��Mˇ\>�3&s�s�U�+Bsu���������9�Hax����*`�3�aD��Ŏ
7t/!��k���8z��v2��h��l���mڑ�]zV7�������9P�7�9w��kƛO�6�,����OI�e{��&r��[��a'�']�وIѸf��5A2�n����!��߽5��F��&�k���&�0�l��>$���J��|�_��X��S2iȋ��yy��Ͱ��Z���K�U3�<�/��:�,����y/WM�B�I(�#OvX�}� 㹗��t���/H���S��z�@p�;��I��i�G7���q�}�#�L�3��v��C�7��wo"l����Ϸ�7�<{[S*[��ᜋ�(u��	c���ol͉Y��" �/��, �j3%3�>���W�P{}�0"�����7IY\����#a�= 3�M*��o>!oc�]�)�Z�{��U]��a%�x�$F]����O��9�6Q<@��0b>��'�gu����T0!�@9cJ/#Ղ"���1H#ǐ�ծ\n����T"��s �����!�����=u��I�N ����o���a��l�Ʌ���u������O�oiu�8H���Q˩��Ny�򀝫�U�	��
�g�Q퀱�P.�R��hS�GW�gDB�h,_]T�½Y(i��{@F��8��t�46�t�꬧Ȍ܃������t��7�	d^��-���eW��x1��/۵����F.�����6��0T�,LL_:�|\�U=
��_�v՘X=�s8j�w�!��'�*��*�t���e(�X������r���x�̚4Б�	Q�������!~a(+{��\Ư<�4�Q���`��"�[?�/n�%�l���O!s{z�B�у���NMO�%!�X?;��Kl�B5�h�����{&�F+r�wIk�����&`wL#���$�Իh�`N���@%�&��?"�!d6�����Ї��D��6W��3P�`j���0q�c9����h��ZRr�=Qnu^L���S�t|1T�].4z������}�q��|�#�\�������vC��~K��"V,�0k�ver|?lŝش[C��ߖ�g:<���z��ë�i7 �=_�ɴ���f��,��	�v�<6IX���ʕ
�i�Wv�ok��p�n�.cnmr�9���1��A҉��]k�=H��3��jԷ�EE���o9yb���Y�5$@\�� ��򌦋J��vL;+�S�ʪ��kk}���fJ}�)�,���_i��P��#���<.��W,�N��ޖ�Ϯ�<��?:�pH�Ai la�,�0;�nR��9����X�����BUˀ��e�?���ι��D�K��bA�����	y�B�Y�`�S&�_�j+~,�rB�*cB�b)�,��	>��<�t�R��~���PP.\^FVY%�@��/���1!E<ĤI�� �2H���rmږ,�~fn��]�+b7��4>GX���}�i�������3fn�R����Y���ف�������%IP>����w��f�Fܟj�q�`w5:�&{�%�^h�r,g�T�tr�>��"V4,�~I��������
��<*a�r�m���P9��:��q��	�|�@�t�?�[\ZY�E�?�̨������;�t�ďhVP��w%�S�����//$vE��ʲ��8	X"9	&�@�&� !��1�d�zt?>��>���@n�@N��{��
I���+į���XM]_�y��?�Qy���j���1��T0��r(E��������p��y*�@��	�Zf��_'���>���ST�Q|Ī�����`�ک�)gC]���<���E��Ma)
�|@W����i�`��]�o�HQK���_���՞|z��R)Ëw���'}��MBx�ђ��Hn�4�q�B�~���ƍL6�y����d�����1��U{	A��EC~廩a\F�Bg&KƥCD���e0�����ρ���)�b&i]٨�� `��x�î���rR�בq��is�������'�d8�e[� Uzw'���L��e8n�V�/��Pۛ�|�?��}7�!#BB�!f$���Y��6U�?��ɜ��ګ�áKp����1��;pf��.�4�f߬�&�,.�I�4}B=����w�0��I̞�Ri�>K�V�'1�z-���$�l;��U�;]���"wt�;=�P�+ra��j-��'OV	�
9�H�9�}'^ �Թz� �ͼ�D>q����	���!w7S�����v�д"@��)S�HF��w{kj�G`6Mt� �Gyh�9S{�]!rD5�8�`UR�SeU��v-	)��Ҁ����h��u[�7�Ӡ���J;�p�g�H�!�g�*��߿K��d9�_E� ��G�Br�����bS��dk��"���ؙ������Ã����c��ޚT����9\�����Z�n�W��KHJ�5ic�kO)��O����� iH&N⭽����I�}���iD�K�e�=&/��A������x�~=d��P���L�ga&���~j�^N�d%��0,��@1`�
��<�)���4��������'eUNS���F��m$�U��U��2
 Fy�L�>/�l��CN� O���P�G�]�Ve�&���dI��M�%���Q=��W	*���
������.�x�|��^�1
�q|��Cl٩�TN�R׃7�����Q�'p~Pv�T��U��7� `�g�=8"F��|�;s���ف���Κ5u��γ�s>j�aN���{?�ݙCܻ?�N��*��X�@cy�L�=��,���<�����ء�03��W��������I�N3
�!��D�JNg�~׬��c�j��(���Q�(�?;~�ܶ�B��s|(�����eh*�ͭ����sb�ߓ��r���a(��7X�&����l���ĩ�5�gR�U3�>w�'/�FW��eV�2!�;��H����u��?T&<P
8�χ&��Me�|
���1��k�<7>@J�|����M���KSN��R=*C�}��"40$��z5ED���	�����6䍢_3K�-Kgs�.^�X�c�N&
�rMk��LS���V��c,8<�sl �Y|5\��������g���C�t+7��k�)
J��&ذ�[�"���LOM���x!�Xċ���?Lk�p6�.��)��@��� �a���������*	 gȓzm��^�߮k�W{�0�B��wʴF��N9ryW�O�,�V���a�;�9z����Gf�Q"�g�:��˻n�
GRh���L�,c��Zb�oB]^��u�F��x��c��.����Y7�U�{�ߦ���?���/���Ḳ
����/9�{�!�f�Vq���I�K_9�]��%��08�y{�-;�����PD'-��K������/�QĀ���6a]2�ʣ�r/J���˭ّ��(|��7O�������=o���Q$�_�(�*���F�ڬ�C���{��wv�	)�?�A~�WSA��O��4]S��j�IB�{XD�������	j�_w�o��K�YV�~�lfqǇ&��O�XX�B��	A\ȧF]��.o�8����*h+��s}�=�0�/�t�3��_4�(V1Z@�ūQr�8Z���(�9e;{��K=]�?�g�����L		�r)m��%3�괌��6���O7�
S���rîb��р$F�ځZLP���K�ꋜ����������� �B�
�p�M�h�����5��P=�~�W��	���X��h�����>M��� �1��w���I��x������#�'_�����j-ZC)BG��b� &�l�Ɋ�p�Ƴ��+[���S��4z��scSRTGGw���+���Sv���L��`��IoK����;b�u�L���	Tg��b�wS׉1�m��RB?%�@ߚ�����ob���ۦ�\r�����<>jꦹ�!L=�7{&�ge��F80���2�	�����_Gax�J&N������ �2��U�Z���D��z-/Od�pB���,��B�ĕ�Kbm���x�y�Z���a4���UVh��P2�[��%dR�|����֫�r>�a'�>g�);�;��"U�:e5wN �Sv衣�9���И���a�6�h
�ҲN��a�؄R��X��6��d;6��j�IJPB4$3F�7c�g�&�����B�H=���n�PZ(���C��]�wچ���{�(g��5]��/���������c�#H��P��B�}�l��ӿo�լ�)�:h��M��ϐm_��P�c>r�x�_��$�>[̻����d����%�X5i��(ې$4����2Rw����@p��K���|��v�v���}^Ӷ!pE47?��b�(!2��$�w���8�-y	E���k[܌?�F�̏������ /d+����E׎#��(�YF�Q�;bGz�4/m�R�w�W-Ԧ��M2�it"�{�#�,u�)qS6qS��}��n���h1��/��؀�����ĔQvt9�Y��MN��'/��W��=@�X�o���k_jN�E �s5W���e��9$�9�W@G�"���h^�c��w[��C(B�i�uk�I+�j_�vl�s�W��Z�����:E2S��u$��?�$����.B?Ҋ�IXlk7��w@Dڧ�cL�Q��(#���@O�����������f�N앎R��XEa��z-���4�j��������_"�̸B6}r8�1us	怹�]�Ltnv�����\�b[>=cG��@��cщkx�dSW�(2�s�<�:�A�$?%!�C�Bip%\�]H���2��/��������o%����D{[�42�i��#��K����ea�]���b6+?rO�Q�ƨ���'�{߷��_�-�d�A.�r���V�rI��ؤ\V?�M��+����H��Vr��0��!E���k��Ko�s��7w7�
�U�6���5U`�KU��^�{ܣ��iH?x��)a�\s� y� ㊒x1[�u���g�	��S�iH Uv{�_�Z��=���v:�3���D�
��V�p%*���%E�M'����^�ױ��M�v�C�
��+s�}��f0K���^ϣ$!	%q�<���B�P��	Q�F�߿e�����_6&�� �edυ?�cM}�"���=�O����`��06�J~�����\�8�,�48Ϳ�+���B}��}����ؒ�@=M'�$Һ��	�dpb`�&])�c�h%�[1�Ѣ�c�v�r�8�&���`��}��ḅ���	�-xM{4��KLɘ%WW��g��-�{�l�r�04[��K���d�o��;��8�\�!79�Gq���#������wR3�5��kpb�颖.�s8�~G7��k<�g��M�:��n����_��r		=��p�-楪�*f�ZDF�
�͟�C��s�ϬZ�X;�fVƍ��� ��7�E�/PK0�_[15�zs3XN��O�%��Y��=��S��w6e�"�DI������4%-��%�h�]�40��ԓ��H��4��۾@P�xD�\�F2ED�`%Ba�A���-��i��h%MJ
@�$�-�5�ċ�L	�u�ʨ�/�E�Bt��l�$^�^�����w�����ݣk�Xv�j�M?���_�dM��P#�Y)���?Ӵ^��J�;b�)��\��&f�1�:I���t6����:���	%Z��W3S֢M�rg}����]4)%�H�b�t�����東.		(�&���>�i��rx�������U����5j����؁��JQm3�
��
�=D�����`�q6_��'�P�+�o�:�Y���Sv�9��E�˟��s��k��ՍΥU�L�Ϟֹ;*���f&�vgs�L��~�5Nb�p3E��\.�a�u�����:*S넯f3���kԍ9�]���Ab����;m�X�4;pB��M��,K�lf��%����Y=h���n��U* ���R���_�[���* ՠ���h/;��y�C��[��^�AJ��Դ�T�\p1C�i)���d�Z@����_�r�M���>���i\�H����fm����u�+R�����m�=X=j�i���|��[�!Y#���76 W��?�����<���w7�3M�AFm�C�Q�j�-f�A�-�u�/����릫c��_$��+z��G��NkX�bƏ?5��$+���0Xj�wz��I�di�����_�߈����l��h0o��z��
���d���w�EHے'� �2@�^g��T�>��@���3W��,��.�6�ݶ�:�,rY�"-+@/\y"$��ȐZ��\;��_�\)����>���� �Md���{8���n�2����_�	m�w��-�M�VED�����cA�<ܑi�=����#N^i�?� �ě]U>�L�Q��h/��`���Mk���p|Ih��'c��a��n�锡�,�&y�Q�J>�0����:P�en⸇�wCes��Ƭe(�z�z'A#D:����x2I~��$�n�`����D�<�;��w� ���&��M�og�J(_-���U�$�`�'ȁ<ҋ���ߞ1N����y���g��2������3�����-#���?8�<��ѿ��Z�>o���c����j']�{7 �1�~�����{*cZ�{47����H���`5^G��,�&����}%fNO����0�4�f8p��s	'�C�;[�ӟSAw�m~S��J���_�[Ƀ����ī݆>�3Dt��^T��w8�{��y�݄�Rk�:�E�_�C6�|H�n�(S'V��ܖJۉ��������F׋�?�_�L;Kk���_/ ������©��f�2�3Иc޻zd�S�[��9G k��[�>aer�k�w#L�E���˕|2e?�ta3
>����g�A��4HQc�N"��
O����[ƴS���v{���'_5���wϘ�~��l������R1 ,�
Q���2�'�Q"���B�_�?2l%�����3=0�)bQ3����h�Zk>'��5w)Z��㊮��VI[�QK'��ZXulђ��8&��VUp����x�m�`�
.�z��پ#������R\ʻl���b'�s����gs=�ް�׸Q~C��ɦ��C+,ˮ���(<���������eD���4��;CJ4�O�,��K��Ǫ�ΫFƛ��#!�g�%06���i�^�н�3���y8����l�T�堼�QU���SJr��ZB�YBJ����pʧ��\>��i���;�h��+�ܶ��2�(wDNm�y�z|�Q䗈�&.�Qv�d0�1���h`�Y������@Q0'�w��zv��n�� �s2"B����A���7UBR�g<�������ʣiY��Vr8#ch3n��tv��>�=�&K{$���/]����]��P"�tR��W��;oO
���7_k���1R ���m�<�����4I�zNY�r�l�rxi�xf��G�/e��O͡�q�fj9��0�R֕�ܶj���[���MX�v�	)��8��f��͆�
�^!���S��w'�ċ|�,l���?k�n�vkxp���㐘���'$�g!B��)�������m�m�;����^�:��{U�qp�MKYp�y2(vh��*i#s�bʡEJ�a�/�}��FLB����52����lR�'��ʐ�O��>|^I��뭭$џ[�^A���6%��r����C�,�9c�(�ׅeu���J�}]B0���X���nf�aA6�'�j�F���V����9��a,��JK��Q����7+�����΃1u��d����dt�2]�M:��_t��zHfֲo��r@'4�����b`�((s3�\��>����yI)���>�Ө#�c�~�_�����������@yRڙn�u(!EaŚF�ed�Ĵ� ٢ ��n�*�k��pƤ�õ�-�����j������n����ŜF��J�q���2��ؠ�Z�b[���y)k-�ma����#	mW��6�=�!�5R�
8�3s#��:1�����O�XK‰��XY��fs�bpl�x�d?���r_��hu���䭚@�Շˢ��r#c�}�v@��E}8]�o���(��e|
G8��V���x�:{Z�^w�]��w�(ReՆ�6���bTx��V����k��Ŕl�!ߩ%ܻ����}5�#��3��F�ɡ��N-8�En-d���K<�z �ٷ���6$�t}�Of�M�>|Ȗ�1�Q"��qF��Ʃ���ȁ�;[u
.�3��aZ��c�u�}��,\�ջ�WB��Qjj����
~&�B`u�.o}n�#݊�պ�4{-���U�o&)P(�Y�-� <'(L}kv1��0�c?���� �O �4�~�e۞Ĳ\��o%����Y'ݷ�v�AJ��U��?U2?�j���J���P��X��-�.���� 6t�X��ڝɬ��m�:�wZ�
q6	�U��"�/���\�2^b���F	
�2�;�)1��:���H�?QP���)@�I��j��q]TWp�+%΀�=f[O8��m���Q�ΰ�	�w#C+��&�.&cN���N�+�_�d~�~lf��ЊH���{Da�W�8/*��'�C�\��=EK?�7���*�r�ў]�Dř�@6w��	�l���4s�{/2�o�e��p��8E�:��c30�T7�#Ye%B*�9��2�o��U
Ĭ�{�e4�#�����P?ӵ0�/��� ����Y�Q4�c��������l.:<����<�� �j>;\G,^a�9�T����zyκ�N20��V�[J�*=l�#�V�J��U(�P<:4,��c�2d�gO�����\c�r�����i#�#�&�$Q��x���oƁƓI`�� ]�՛K3 B�	��U��ӗ�vN��g��׏�5�����I�d^�8���NNP+M�K�P>���Bd�3�ڈ"ϹKzz�w�=����t�^q��y��d�</;��c���/N����/-cW�-�}3�"9����=����Z�=���/�L�K�����Q�&i�r���ڥ�����ROw�
�S �@���W�b��(�f8��P:��lV�CRB�!Fy��z�U��r��:��J�W[��dd}�������$gӟol�>�Q��&��΃���hն�e�w�!ޡl�×�i����Ae7]'u�H�;��Jz0����z�Z����ƙ�2 ��zD̑���Zp�H�B�,b_�+�M[xc��ʪ?aj<���bvO/G��^9[�,�j�<�Wi�т����P1<�n��!(�_ܩ��qY�����.#��쵚�G���n2U@]@��(�dq;��Ul0P ��(�I�0��xH�@�*�����Y��{�5a�]M�2��^�^� �l�R%ؓbK��j]���Ox||ak����u���oH>IGî�ĝ�ƛ�I�]��wL��ϻp��M�߄b3r#���oB�B}����.c">�"R@E�F�P�dݚ�y�[8�����7�v���E���QL�UZ���w��܄��Rw�������OU��Sg�{���.}���J��d�?&�Wh+�kEA�ݢ-�M��u�E��������nWJoڪ�x�$�/��%��Z#�~p�����\
S�G	�sU��Z?�/z;5>�/�̮"�ѹ��-�qdu���X�&YI�,qz����"nz5�BN�~C|�Cń��ǟ��{9�.`��)
�q�Aȃ���܂��h���j�k��Cò=3�Y�߲��ݪ�j��c��I�7�d*�/�獲�"�9��H�%��Eђn��3r�W�4�<W�|�"1棖W�b%�Q��(����M4���XVW�b6�X.f�x�g�D��w����&FF}�F�HU&%p�q���\H������l�s;����k��5�w�_z����e��Ε5t�?IB�>��2ؿ�	
�H�R<�Nبe�q$!I�2&z������P��^�P��Ic��Z�7���2��i�fL~�b���a�� �M��Vx�@�|E��h~�Nz��^]�16x��g��jb
	Փ���Ε����kXs���4����0�sޙF��󬈕�����Z�*Os��j��]���%mƆ���WCPq�a�T�R����J�����\�s*��r0��w<~�o�����j��E�f��_]��|�����C2��s�8XX@�i_�Bw���Y��#�2V���]^�5`��龰�4
B떥o��%�Y��Э��Qux��p�Љ�5���RZ�Y�˻L�B�n4p1�P� �qQ�p/Tc�x��u�ty�r��^��mؼ�]Uz��|�����
ǹhM���9�����-q�t��)+�;ƨ�3����)K�jN=%f���wj���	�<�s�I74�r�⒫cj?`����$�o�Vº�L��e������{U$>H���?�7	dy�j��X�^R'��T~���FR{O��H��%�WΚS��y���~8J�������k���E�+XKN,���p�ú��#cY���N���*��Q��ڔG�f��Բ�>��j�/}EZ��T�$w��O�/�mu�"�1<�;�v���L]FF;x~��eg E����,�;��K�,��ʭ��iP��F07�IRO��$6X��+��z�E�hq)�i']�Gw-Xn?�|����ڇ�����ۃ/�VE��^�>�x���IN+��X�2�1�����HJ?ދ��Bs߼�VWJx���U��̷�d����uX���VP�1o��r�ŏƉS{	�����>kk��b|Ool
�EL�
9�'�V��F��:��?#qX\S�ξ�,�B}��w�"���O�v���i9�W
�A��`(�]��>�t4W?a��cB7t^��ôv�/i���C�7�-�3�|@�����>��ٵ:}���(gQ^�2K�m~���G|궖���S>Iܰ(���c 7�< F�e�@@3m^����,���p�_b(�j;�:�%�N���^=�����^���_SX�I�S��u������-�<k�11wY\-���dҨ��0?����ś�	F�Ռ�A���ىgL�M��I�3'm�r���y��>��}��[8�����ׯ�CI�ث�S�)Qa�����/����}���H�4ÚF@"�&�y�gd��k����g\Z�h��$_���7m�Z{G]_��7|���g�w��5t7~p�Zρou�%��i��<��`��o����^;8n2n��K�_����Ƀj�Уr#�]��q��v:<i���7���ߐJ���������f�M�á���A����U��ˎϟ�<n̓���-��Y����Bq�;��P$S�g�g4 ���=�G{.t��e�֙�W���W��+3bJ@���af��^�̓&=���@ǽ�}�w����5I�:x�ks���`̔Ѻ��2�a���S����94G��+�]}�ƛ�<����A��s�T]�p2i���`��3��;5،����VJ��c �V�=Y����'��:pJ�o�pq�}�D��&2V�~�����?�`j<�����M�N��]o������s�� �Ն��؁�k ���xd-�A�#�;�e��o6~o� �k>�1t�C��^M�M��$�ϳ�+�ަ7�'�L���U}l�q�zO���u,�	y�O�;0�p�ռX�i�?�{��eM��ҍK�D�w"hJA��ʾa�)����Rt�jC��s�k�j۞�mm�սQ�R4��.2Om��x��yc�ϻ9q�K��`<�	/+��67Bb�Ĳ�Л�c����A��ur���3�f�QI��B�E}����=�fA,֭g�W0j������j$Bl}�5�s���-K��[`<Ў?���.�5�q
ǱB6}̯���sq�H�%"���q���`&1L&/~��A;�`�b^��e�\\9�`��������<X���җ��<�H��'4��q�&���ʹ4�^{�e�1o�ߣ(=�y��� ��å,�JJ���J(��M_pN��Ϲ����p����m��:��4�]�5�����S�z�`ϣeQ�Bf�+W�4�̜��k
�Z+:��&��O<kc�T�'����<�J�j���g٬O`��l��k̼x2�J�#3g��y����D��#��3��!3��_#����p���+'������m����k5�sj5%g��36�Nֽ��Sxe����=��HČ� Ȇ����pd=9HFr�(�e��d���x�QW�6�0e�3v�&ϸ��Q��}�i�����qSI��'��e��������R��9��nfo���wI������6�9��|۵� rz��UJ>i$i;!!C�c`	F$�a� �Z��P)��Z��7�{�m��ރ}�T�覈ih�BF��r7����FF½C��]���j�(�|J��� Y�%Dk�)�u�Hp��.�b���T%5~���/�=cɗOT���).=�cJ*L;kZ]F1��O�b�aRkb���VS��8f�!��vM�{����C��jL��������ș�?��S%�0���/�ۺ�E��r�>�4����s9�R�E�|b^�|t���؅�O���r�h��mt7�N�I�])Y%��tM�t�h�����A�@Q޲�3عx$5I����㸬������5�7ym��{�w�B~n5��l�u�о�{i�=��^i^��%Do��S�<���(��#�#7]�"�O�������HB'=��#�b떱���}�����y�s~�0U�����X�S񦀚���`ЪGn�W��
HC����!{J�b!�a/ֱ�ۓҨ*��l�>ci��~�v��I�����G,�j|�t��%g�A��q�=<F^JR�	 ���f4:��SZ+vY��	?�����y��=�Pbx(E(�{{Gk\j�^J�-�^�q�j��؜k
ř�����������s��]V#:d.�|"�^jF�b	�[�CM�w���V�o�6�����~u��|%�P^� Y/���F��j�#��*@RK����-�	�9�cJR
s�e�����x�/�ևB�4�� ���:v>�B@���T
:=��|��v뉾p ŏ�M��L�$�c���|b�q�N��-�3L/���r����l��l��*���9�:���(��r��"��v�4�C�U
TTYah��*?J�Q���X݇��L�q��P��D��ϗ�&�C%)��q4{��� {����Q��{u����x��Y'������U��>2~�����I��>b�3�y��F�Ig<o�gѺ����I�$�ʥ'���6�+�o�2�M�;0x����js�ڼ���׫2P�zb�`wy��HޖՅN��4 yz=�R<��>:<��"�I�((�A�O�� �y%J��Ş��(���5����y�Qy��zP�r(q*� (�vQ��C��?S������׆4���u�=���|����7��0oJ�"�O�N���z`�V�"��~w��k����� ���ާ�[JB:E��K�;��AZ�\J��^B:W�ARR��᫟���g�;w��{�3w�L�~�G�6�d�0̽8�䄉ls/o�݌�щ���R.!J�������ߟ��|>Jg��I���>�1��;���S�A]s+I��Zj��w��EGJ����O��C��`w��Ż5Cx~��������Ѳ���!�>�ap�=�u@)yQ�H0��|� �'(��/���U\�]��l�R���$���u�gzd1����(UٜjGK;`E[����
��Sb̵n�x��C�:l���r�Ap0�����5!�.��wN��a>��w�F18���w��#�ﺑ������@YM��'/����[\thQ���_�C�̖�ЖZU<0+қ�-��K{�A�lѬu�p�5A��[қ7��2�n��犒g�~�� UW���I{+���@��C�-��&ذ�e�g��lXC�#�&Zһ���*�Q��,��.>聫:x�t��z\-��h~8d�v�X��?7�/�!~xJ�4���GB�a�6�6N-(^�xAٕ�w���+*m�OXk���=B���YO�;Q/z:���䪉+u�3�գ� ����Ib@�_�3��t2.�N/�4Et���"h�s��d�"F @p�����x]�L���{�P�`}$
6J�݊��,�՝��H����q�3�Ц������"fʦ� ��\#&(}v�7gMS��'v�Sy�1򫅬��׋E��S����=�m�hR�W���������`LlI��C�z�:�R�c.��ܾY«����4|�5���P#l�_��ϛ��
�ez��Ɲ�λ�C�*��tG��l�7:M-ED 0�m���V?�n������RԳ2Z��DM|�ڲ~p�w@󬂿5K_%��
�v��[���l	��륏&㗉ۤ�?�4?B��AA[��熑���ij=�\A'�,�@����г ^i��)���s��aĨ��.�j�^�p�u�mL�.�Xs�o(>����ꅺM��i�R�z\Q��|^���f�9�usj��\Mo���/:[Z���p��i���]��-�Shp�x3��'AX��~8�ٞ,١Fp]�L�����	�I���;'tY�~� ;T"�:��ᵷ!}`6�ou��j���$yo�e�wY�6R_Q.����?lm:���]��{5�t�A�Y[K�[���?m-��ӣ�-��ӏ�R[H�νg�^k%��-bF%����"AG��mfڊ���h��r��	3�+8u'f7�^�;�ß�1T�$��\@��jE����&�[��H�rI�mv�\Ǽ�̚(���z�t�̮L��=X����䀙,,��sk�Z��eX��Z�L 3ʖ	��{g�r;� U�J ����ٱ�,CL$ִ4��z���[E�D���{f�T,��%����\�+��J{�>+�����XA�QO�����~�)g��k�\�ԙ�%O��aoY��IvTAԕ��7y�.E��8�4��힪Źn~�w�p6�|�8%vk�6vG9E�#�}�}S�]�&U�3�u����&d{ӆ�m$�r�x��
��L�rj_eā��Y����M����D/�媃/4��$.����QU�Mp���:2O�q�E�np������"����Ill�=�@!����xrlXw�Oі�h��q�q@�������+�7�ao">Yp�-Mj~�I���I�u�e�%QFf�9VMQ��ޒw�Ô��=���|�M �@�R��Fo��:vN�7p�$�E�&���De9Lz�\�W�0��jS��R�r�+ûT��让��}~ؤ�� }� i��F�� �E��*D�*8�SY*u9&�y��g`�(���v�>sD�u��F���̖a\-��<+���0!֔&5N��J�.�OpV@� ��{ѝ�������(@�b�E1$�S�tvw��E���_~m���㇟?�}F�������{Zs��wK�Zd�����D��|x��[�B�Ҵl�D�Z\�>�E���
R��!�-��Y�K�v6�W����*��xR#��_��3}�.T�͏h�-1v�B�ٶH���O��|^gɺ/�r���ۡ�(������?�C]�䠆�N�
^R�uۤ��6�A�wn/�R�w�'�{#u��"�~"�s�f������FrD~��nϨ�V��W��g7�Ҧ�?�-#���UV�$��(j�eR�Q�ܻ���O*v��T��W%5���es7�&�.�0���Eu��n��6v��q/�Q���9뼛\��/�OO�F�^�t��A�=w�|�S���x,�n��K���~������3J����^��	�d���ۉ;���,�μ?���8)�#ϬV�:(dƃ9�'�dES�V���h��"Gܒ���S,�1��*[��]@ĵƎ��ך��  b=j�S����fe<1�N�S��i�����@���q3$���p���^ȖQ�1nMNL�`ηc��C_-�5@�S�ە�W�1�UL���~���*�������S&��;Eցl�5����W��U���Y$A6y$�R[c�Y�0Jqa��t�����,qɂ���}�ܸ��sV� �ɦ�6����;P����+�=[^i8�{d���v!��8�s�SAV�z��4��a��~$����-�7�����:��Ø�<o���6�����NH�}ElG�i�쎑(�#����-sr��`s��]e�֬���p��Œ�u��zAq~Q���9����b�ou�`_�s�=fd,cJ$
����!������R~��f�`�1���m�A�$9\�ޝGW���|3����2W� W_w=A`�{WzKQ;�B�B��~����7V�[)�l����j��~��#�Mir
�&�o�K�����~K���PG������5{�%	#Y�$�Ӄ��v��3~X�B� �w�(��wsTbO(�T)�|7���z��p�|9���4 и;������o�7V����V���e��"͑�x�K�u�ݔ��Y�_1Q��)�!}8��f"F��vl�HG)e���Z�[����(Ã���0�Y	���Ir������(o{�ˈ� ���X:��?��[|���7s��$���Q��n�Pd��I�]T���I�2��F�|	�M��,��@���:���������[q��x[�I	��i�/v����'<5݆�Z?i�m��Ct�.:�s�Gfa$��rtt���ywSD��H6)�Z���]N���D��������Q)�8�Ǯ�c�sb�q��d���;|ۇ�z�Km	.���D}�}�%�V��`��r8�f��$j����PO���h��q#��MK  �啁�l>�ӆ�C��|�XOU�us����w]�ma*}��2�ژ�E-�G���݅ٚ��Y�t�=��:���y��J�R)n��=vp���n��?>��|��1{d�����$~��q�3O���Kmd��uq�+|�&�4:������jiqk���uKH�yW��h%�0x�hYBq��N����f�n��>�9��_��,�,���?��o�P΂NMn1��9Ճ,�;}�\�"��@bp�����\ܗ�^���˶�8K5���|0��M֞��	�������pr(K和<BGh�q�(5Q�YCd~a�]�,�ŀ���}��g� � #O�C~�t��=!���/������<�=�E�: p��|���Q���6>\��78����lU����IJ�#����Y��"�-<T��f�L8d���L��ĉ�;��>0��e�啛��Iշ_ߕ�m����$�"�$��Y���ei���<ώg=Pl'A�g�Y.�U4m4���#$N�K��7W�W�e�x������چM��;c�HsgKb.�Y�6���.��f�� 1����OPr�]�0ֹXRm��IGmRŎǞ�5�D���1�-[;Ǧa���t�A�[�{�t�8�w��\�I����P��HM��d�o�Ţ+W��&Vm#�`WgK�JY��q�Þ����oT5���0�r(3y��Qlv�R��m�?8�߮�<�������5e�������M�+���U�6�D|���s�� [��t��˫���,n���V���Dx�73�W���Z��T�:�it��}O����3��ч�v~_]����wC$K�1��� �����V-RJ�zԋ���p���2��`�/V^��x��.�
{-�Z0�;L?�!0���ɼ5�ϪȈ�WVb��(���gu:En`�
�_>���A����pD�ArFy����<+_X0�h&ה��͇RT��/^Gm���{�]rr���*b����"M��wD�G��/U��6������6{�C% iMJ_���@�i����C��j���ݗ������ڦ�����ܻf��ψ%�0]W����5ިt��X�uK\��۶�����%�JYW�A�E��[N�W�� �pǦ�_k��o�۩�/��'=Ā1�Α>�t�?���F�0�{�x��9٥Ƈ���~7֊���`31����z}Y�R=�������9�ʴo9(9~x��Z�ꝲ�~W���9B(ӹx���Y�� �X�пYt�tAn!�m�����"µ�E�4m�0A��ō�f�^gY�/��za˒m���Z��a��{5�hdoEt�˖�W*��n:Y����8�]j��ݥ,�������c��0�*Bpӭ��?uY�m+ 'dϥ :s�q�f���(���!�qC��;�V��9����.(�)�[�E����..���>��;���~�|[�9b,qs��/�W6��n��u!\k������h�9���^'B�m����t��W�TN����c�>�cE��[��h/e}Y�ɋ5-Dƽ"�.�w�-r�~���ο�;��N�����uV�u�W.Ew�/��$��� s�TR���F7I���ħ�8*�*��>�fi�j�O/��bq����]�~o���n?��~ޑ��j��=�s�U����΄�>~����y�~�>a!Y٦DOǏ�ebP�VZlu)u�v�/'M���~h]�J �"y�(� d��u^b�*����%O�+�o"�)j����ƃ&�J��|e��j��zL����.H0�NVZ'V�,FV<�*-�}��%��¾XҔw�(��n�$+��,@�;�o Aʒ�0!�Y��e -;F�%�r�e�v��p �x�}�G��>�=�t�$�Bm�����Q��g88f1!wF���E��@cI�7��$L	�c�,G�(.2U��JK�}�&[�y뭊�bF�,�=����ieT���\�n��K�+�����=���1�;�w&A�K�ʢ�d�ϼ+�y˛�q�5�l�{{X|.���=���N�C���?������9�O�ؘ��F��P�,�1m�H���7|C��'���������� ���Rk ��*~-���r�.�	/������E�z������J��k��)Gf\p��m�s7�T��?l9U�v���Mj��iB[R�(�KX)~���J̒���7�g����/�i�۰i�	��&+�q۩�]nD��|a�<>�5�m�"��J�����)��#�Yvt}�a�,��1_����RN�$�Bc�JiRO�w��R�%�^)� �˥+§U��X�
�a���_����n�\~m�wkV��if$�h���G��J�w�y
����x�lY��ُ3�P4�4����p�}鶑���kv��B/�Z�rs�[�nM5���<-�Z�U$���Z
a��Qέ�DB=�&�ߒ��Z�7��P��d�9V��R�T�bM�T<�Z�%Z~���lt���BNZ�@o���A�.�n��	I�|l
��!�j���f��j�dz	�gzg�˟l3.�OT���@�?�gL��X�eL/'҅b�_m6�a���$Sg��U�l�铝�8�֠snΤ��a��\����UA�(�6��ɀ�]��/G��"��ޛc[4�z���w�)�@���&-N��g�n9�=;󠨲C�@e�b�R��:���d$����!��BD6z�ұ���{����U��n��ˮ�;.s��X�ZIϵ�<���3ܘ�П���d^��79gNC% c��j�QD���`,)�5S�-  ;�hˆna���n�?�x76��5�j�+��@���^���(�JO'nzD|h�Q��Ӈ���XE9����n�Bt̮/Ҩ����ο���+'�Q`@�Aސ�n��{����.j�x��F��
�77F����.>�+��KzC+�y�=렶�cf��Z ����0�����'��9!}u�SA�W�9QeT�QrJ��Tz�	^r�$�՝+.pt�5�����FP�f���Xb�Nm��4<���k]@t5s?ѴBxn�i�o�C�OoȾ���/ G��.��Im��/L����B��Ӝ���(ݛG�j�B���J	�qV�qq��ţC�cf"@"����?�����g=+��Z �f���ݱ;��|��fuU=�oٷkya��DWZgT��jFz��_�O0��R���:u�)�#Д_Q��2�ʛ��Ķ� BٕU�v�k��,Mɤ�+t���� �G'z������!��-GF�e�׊^��mf*��h�D�Q윂W�y�-�2��$u��z^�pf�R7գ�/N�I���-M����f�/�@�f�%���;��O�&��ZZ7}�/ݪ�y�;ͬ��=��1#���nt���􅢚�up'��/��+�e��:�v[l�L�<�н�;�}l�{�R�JTݚ7lWNnX�uv;�3��kV�kٽ���_ui vϖ?��M�A�QX0ʂ����	�F�@8|����A+���-tT��1^��
��+6:���_��]i���vj�3���}��W��@��D��2���k�Hb��+�w�O�EN���>��[u�+�T�B�
�k��,`0b?¾�Q��yQ�+ܭ���2�t�΂�x�Ғ�Fg�Y�h<Q� [�+��#���+d��\H/<il�_e�M��*zWe��%M��Y���Qc:�K�y�� �A�A�i-���=�ԋ���T�L�C�2u!hr`���{��Z}6@��*#n��;ԭ�&Z��=�t��l�4�+m�}�FD�R����<�X�Sv ��ݨ�:K��O��]�/�	���M�n��_�0��t��z{�����<td��<�}s�ПPP��u�\f#T��c�P�^��w!޺�_�y՜z�d��������>�c�L2{�V5��5�$(���gL/ �Q�)�𬧋w��1 T�5�r���-���]h�+�0@���Ш+d!]����=���*"��6]�~_�O��7�ܝ*����ZRZ�Q�W\�̞������J��7�����[8M�B��JE�A�G�C���F�é��Ǘjxtkw���_��f�ߕ{ƾ�_�U�w	s������.eu�����4�3�q�fO�����S@jI`�!{�^o���ݜ��vN���h���;��4�KCg�R���)�TT�o��(U"h� 
��Ӳ��|��s=��x*�i2�ֹͫ��4�]��뺯�W.B�H?���o4|��m��F��q-���Q`�������&� $E��'β�^7�֥d�:��G��ܹߢ�2Ćy�Tg9g��c����~r0;�}_#W��q�����ٱ�W}�x9E��3�d��l�^��j$-��� Ice(�;��}vi�=ª��4�:�(��"f���7]�eqW�B��Rth�a=U8A����4.�������ѻl�o�ed�|����m7�<����J&��)',����.��CM�uz��=�a�6�������	���L�/#;���rP|x˷�j�׻���O�O���v�hl��0���+fNbi�
�|ۆ�m�z���|�9��KXY��ʾT�2����g����?��/[��"�;j�-G�j �)I�� G��:�
�rMG���Q{�m���uko���$'���\ʷ��-/��~W*y���j�?ON#�m��J)���7�\��6�|)��[z��i> hoz����-��s<�)��M�Y7���׵�������,���~\�^�FG4���� b�yX#n�ͧ�~�(nja���}��y��b�3�ҹ7+���ڥ����"�a�w�#�xd�V�����̙�I����ù�<�-m����{#� ��~��	��\��@���"� �mi�:iS�F!���K���I-�o��4��L��x����$0+�s��70ɀ�;y�g���8�<��q�r�o�J?-��c`$?���00�~Qh8������w�w�1��Ol�� W�׳�t9�3z�7GB��]���L��=�b�=b^KU"	O��^�)��"c4�#n���f�4��a�%9���_���^���3˳��0��2]6��L:�݁���lt�tw��߇��;h�����x�/$VA�g�瑳�<Y95�g�/�+l~G�^�cz�H��������z|MxM _�K
C
�fUXF�j��jR�/��&�l�@��<*�#��>q�P��]��)�_B�#��B��|�~L���|xoa2�Y^���9�c�� �^ sd-�W
-�e)ܗe���΋�A�8M��9e�0� "
�����Q2Y�V�z �)<\
�U������@�x�����ͤ
l��s�D�7ν�x��
}�S�}x�T.#Y�@��n��0|���Ī������o�c�ૄ�w��i��D��
�@��X�5y�����r��q��W�J5`�(z�;i��]����Q,��0��Q����XLda���zk�{a����j���\mdl�=Q,�h�Tj`�d%p{i&t�)�+'7.��
�� K��=_ߵ�	3f�3��n+5�c���<��� �l�ܛ�>��7�:�l�œ>O����׼�`4M�>�N�X6�U�z��ź�a1���ibs@ڪ�}��}L�^�y��K$�N����ȯ��pd������b����s��R[*+x~7����r�iT�1
0[\���+�,�=�X)����f��Z�,l��0H����gx�ޝ����TO��+�B��?�z��a���o�1O"�lX$/&=˷T�K�B_�z2���D ���%�x;]����tc�]	��m�o�\R3�z�@�\�_��YfO��[P�@�������[��~y;�`8��z{�=/�0��̥ƘÜZ�6u�@P��|l��s����4_*.�hf ^��׻3a���e�s-H~�"�ԫ���ܨ��<������'�O6�M
���	��ZY��
��)��n�gg����VX<�x�xP� �Ue�O/���v�����H ;3�\���l2�мa�jv�Ώx�Z��m�� �����cI�q۹P�4�+��T�~4R�����>���Ď��c�K=��@��V|:L&v���{�_��/C�,ڕ�AV�(���V'�ºl�~%���5�d�#'����?�����}'Ymɘm����N2&��5���N�9��r�Z�K�Y���嘞\r����^���&�U�L*{�1�h0� �z�PX�w�f�PR�L��Ԥa�\����x��T�$�F���{��j����=a��� d#Z��ƨFI�B�y��u6��`�q��*ԞV��L㹔:�A{��A��B��($am������ο��m�`��+y��*W2S����gk�s ��Ԙǋ�$ӫ��5N%~����U��8͢�kI�kT!7�^!.�{^+���s� a���*G�e��Q�F'�Õr�ob���'I��o}�KF�r��<���|Zz-����	�$�+_B�n����W�qT'���LK6��k�T�-�K��g˛�N截0�j����rk�x��:N�]���h-�i�/f��{���߶��ּU�gO��ߣ[�� ��md��-�V��9�=��s��5��.�UU�� ��:���1��ߠ�
�E�.wn����(�Τ��/�>��Oe%�+��s"��N2�=cQ�{v�S�5�X��9�o>�<×��b��ͽ�h�b��ٻ�L�d�dک�ﵟ��eW|����pq-6�-���f[���z�`j���M���W�d"�9H��` �����8���@�����Df�X)���r6�.-oEf������������W�*�����W听�c��}�1z�o��"vv�8PB���/��E�7��M$��0a�����y�}�*��˭K����[Z �f�.wk���k>�^>�'��b��bF����a��o�ܰY���ڄ�7��3���O�G~zȍ�;���{ߍXf��w��d���&w��_E��y�#��.-�3�v1v���'��?��R��^������=W"�t�M���4���޳�\{��{I�ѱ���`�$BCpV��?���(nNԘf�ςph����[^ߔ�ڦ��Xj[c;{$ǹ���C���xs�Iz�K<����K� a���'�P������_�i��)��	Clz'fl��g?�XB��*�r���֮K$�?<`�g��� ��o�4k�@%%���E���?T7�g�q�i����0/@~�~dl}� TFY�@.� �|6���dD�T;"��نF(h�BV�E��}�����:1�_'ؿ�i��� ����3E`�'�����J�� �h�ʯ�!0�GG�g�b��+�x��_��Q�H�RJqɈcA_�C��<���U���!�eq���z��tr�h/���E�$>j�!���#�
�\A�ı�&�e;@��r�^���{��U��`s��@5�Ѵ��[�:�Q�� G~�l�)g�<��עE��q~o}s��������ży�eH)yE�7�z2�j}<�R	+���f�KJ�|���A{�����9<��~��Y6����w�9��#*�$|R�=�����,�䐴��To��Ċ�\�� !'� +!!O�n����rpg|���� ��3ns���h/yOA�9������o�{�"x?>\�|�zP�2�����C�֘�[�;�l6�P�=C���;�,>��}����@�Y���gEB��Т�(Ur2���A��f�	�.#	�8�^�����iE<d�|�?0�l)��Z>��f�$�!�K���أd�EV�;��E��Pr�<�!4�&k:�5f�BO�VP_��SDx=���d�^�\^c���A2��F��<&�L=|&�y�H���>iYӫ�T�d���zU�T�Ppܫ<a�:\N>/��Oi�=��Q�;�W`��[F��>��Z(X?'8�J��K�0�5�$�;���F2j,|$�B6����%��Eϡ.p�g�L{F|HH��"��g�Z��<N�>��CK�����9��+"�G4����5��T$����|?W��W=<�J�w��:0��x�P�he]�t��V�v����)m�?A8�h��{MX��k��p���mU����l���o�Z��ɗ9jy�a��w�5����r����y+�{M��J=�m�rɚϨ�6Df��g��o�
� P�^z�iBt'�e^Z+�F�c�.��NS+l�����I^	S#i�`Lhg�#�D})C��\m:X�I��p�WX�k;[+�R�N��,!.�M�����k���m���/��Fs��pE�}��U2��ρ���N,Q�DR�`Q?Ǡ&Ġ&G�BM�3����+M�#Ɨ,͐"��e�q�MlC��?Ϡ�j�0��m�`�WIc�5`�w�L<2S5���,ẉ��\D�%-��q��y�t�q���a`f�A���R�6��D�`m����+��̊ݱ�Ho�t�&)R/%K�eX�UvV�K4��R�$�:$u (7�ٶk�7�<<�TQ�C�E��r�CƲ�O�������/�܀{���Y��E�vYY�	�2�
�D)łT�<��ӛ�9>��#�Uӂ9H��<1��>dGr�DdBxo�Q#����]&��4�	DCK�#X�J�e��r���e:32�J�.f���]����
s~��:�Lш�j�t��p1;R)?�H�v��8xШ����B�r�@�|�-O� ���hy�o�ZU���Fkޑ�>���.�,a����@�52>r,��x�j�u����<^�e->�h�~d�5Z'ʈ��2{jD��K�0����3F�9Xpq��"m"K2n�f�E<�~�=v����8Z,O�@��3�#_F�Yy�Xs���[`�GE2��HI�����W�$���K4�Ħ%{�E��Ȟ���O�qr�uW��I�z6�M"�{������g�TTU<CE���Nŉ�!��,�X4(��w��H-���
�{�����ԕ��Q3�����܊i��+��;@�RR��}�ȮN��p�|o�J�3�.り�8���Ꞿ������w-���e��H�צ�cy
Zcy�yڥ����S
��K���M��dM�e�o��$l������Fb��Ipp�"Xa�?���FX����\�&�
p$����DGWYQ�eF2�r��as��%��x�vm��-s.�2����WɹP�P(����&�s-}l%�Qt8��3;?�w��ju�7���O�}���Y�d����B�ޱ��|J�)��գj"?�w��}ٔ�Y�*Sx�0-���4cЇ���$:0JJi��}���d_�L�7&U�*�zR[?��%Q�z���)IS�QF�rd��Q�3�.���b�;̇a�}f�H��}���2������&T-2}���M�	�O�x�ae�A�j|�ZϚDNe�ў�M��1���;�o���}���"=�o���T��Ik?S|_X��bj⯲`��1ޏ��Y��%��/QTS2,\%!E(r�����k]8z���?��b���A���@B1�,!=;z-������bP�k=���'z�)�XE)�GaI�����`wJ3���?IZ�|u2F��9l�m(�0�u§q���>�j�S��B�S��|}<�ۼ�J�>��HW	�~�=��M(R�����C�X܎��f�
>u�&�C$�i�6�����}�8��1�1�/�w�bʤ
�5�����X>T�p������_cfXE�#�nD��A�^v�k�n�;F//&����r���y�Y��g���>5`	n�}S2�ǵh�!Uևy(��!��s����*���޶~�'��Ȇc(5J������?72�P�-RkRrZ)**��GןJB��EG\����U���6S�-)����/�Z�1Xgy�o�"?�E���Ǚ�x64Y_�أk��xn��q[����|�m���������<�s-�U���.s8�B��tn��U�;���S%4�X|D�i�!��lZ�o͢R��e���Z�"n�P�MY?l&�gvy9�c9|zR�%OJ�K��Uj�����D/�g�F�� �ǟ��*Ԟw��.s��?�lVcK��za��J�,����a���zT%^�)@�\<�e_2��K��ss�|6*gB��
��r������eܡ؝#���x�ҙ@f�n�	�5ْ�ּQ��5�a��<v7�,I-0�� Lz���XM�}�%
\�jx�d�.&x2���xK~ǵ�t�q�S1���*ӧ�Zf�����b��%�Ů"��S�����	)Qotz	J~��O���_�
���:����T~�5�P>e� ���=U�&Fu| Ak��q����ڛ�e�');>�)��⅝�5��(c��G1죠&Ĩ���bU4[4e^m�+����t���O&&�x���S���^����wz�mñѻi計?|.�m�n~�_/��ę��ei�Yߢ�����9߾�����+X�u���WUb5)7��T/������ޏ�q��
RR��r���_��68Ț�X{niP�����������f�U��Kiz&�$���%9�C�@�ώ�f�b鷡a���M�෈��LH���]5��b�8�G<�}�{9���&a��>G$�/;�0	�U�#Gj��Yѐ����d��4������
��� N��q�f��m%?|T��{N��x��c�C/!|	�|[�Y }�F�X����r���he���!�b�nL��`B�����$2��oU��Pq��p�����,I$���9Mq��=�
ō�P�S���p�nދ�6D����x0�� �h#$�.��`.]|F�z���Y8�T����2X�A��m8Z&����%�?D�_lW�X��)�=�i�� |�(���LW�an1�v	�-�`����"6�OL�=0G�ȇX9c"a(�KY%*��G'V|����C�����{P诽��f�\A�A�*�؁���D�q�ye��B�֭��q���gqdx���(CC)�z9��P�t�@�e��"H��#e�o�	aȗ�xT�"V	�@��G�%ܞ5��x�c��>y��������0��X�%��tt/xY�*�eĀ�B/��Ø`�?�_�"*%bQi�v�u!-��nYjL��
&%��/CM[3p��C&�s�vǩ=׳ͷG������b޿7��|I���f�㟸�)�5V�b1�]S��ߤ|w 3��C{|~A��Sc��8*�t.2����wD��j���eV����S5��ݤx�7�b��t�i?�sg�v'	�I������J�"����눸�m�5�p�����i�[�W�坘h������ġ[@͈�wfB�(п�I{KO�޵R	P���~֊�9��>!윭3�£:F�&�5��1�5�>�YQkJ��6.m��<�}����bn�;ҧiM$	�Z�P�Z����{3�Ġ��@&���4�	��ݥ��IL��ߩk=˘��`�i�t�K��p�F���"Σ��I����}���qY�c��ix�� �52J哽�*9s�1��v����S9���������@D�GJ��i*G�Mt�2�@|�"�d~��P�q�̼�,�d� ��>ݩ�t�NJi�]�I�=�C�2�s"7����!����H��[�1��)��a`ڮ2�rݗP\i���z�5�x^�(��O��P+��[}H��PRuNWc 
T��t������GE%|��l�t�\�p;KY
����(�t\d��y&AD q�U����v�vo\̾I�^���HO�"�Q��Y�Պ����I����+���=��*��B�ؤs9M���a+E�j�7�f�����'��N�|L��]��Ör��yS�.��>�̼��p�Hf�>�͋����L!�Yhs�TC�-o��9|ע��
���#���"j�a`�W���l��AJ��40�ƫIM%���e��K��%�(,k·2-�� B�d50�u����g�i��|�C$*��S�߱��ˀ�ع�U������,�/���R��Ѷ 6F
A8�~��N�B�>�.��;&Բ�4*�\i�:"��Z��$�zz�(�/S����g������?j/����:�F�A.�xF��Ux?R�n�_0^�)���}?�_y�d��Z�t#��a�LF.��푀ԯ�Ƚ�f��	�UXZ��b�B2 bD?%X��{��KF.{��?�^֒�Hpi��2�°1h����B�Pu�?y�M�����$:�NAx�؄1w�v����Y�w2�O3�q�h� ��7�g=�#C4���¥�ΦX���!��?r�L������UQ2O��0�xeY�G�Ѥ��+�_BLu4K�Tn��)����ڳ+�q��������f+@��aD0��? �����C��,QT�&l�����M�IwbL�D���5j����m�� 5��.�1�4�w�z�����|�R�۰R葊v�%&e�ǥ�S���7j�4�SS,̀�ؘ!�0�ad��V,�$;A��$F.�	�N8��a�H){U�qf^&(���e+ҭ�� ���|�53N}�U����]�M�lO�V����0���򪄘��	�l�EdE?c KBt�a��Sq>eL������?���q�����N����3^D�gb0����^����ɋ|�%I��lm�9t�n�K���A����_|��h�1�(d�Ep�3ؔp�ɼ��[�
���E1�����fCMC�����~X����Mo	��Uϗ�Ӌ�n�_W}�%	�LBKA�~0ܼ{"�ԏ�B�]���j�@`D�n|y��l�j��q�?��}��M�
���+�8���䄰2��Nl�k~�)�H�ҵO��"\�Z�;�:ޜ�p��(���6d�;0��L<,�i��ⳙ!)�|�ԙƂhG3��"��;Ͳ��?���>�;��%����Չ�g31	)ɌW��Q��>vj �~e5�.�"�
��ú�n��#t���T�0娏���ú��S�K�C@����%�����&U��j)οi��|��Y��Afo-Wz<�s����h;;H�l'xͷE����U==�M�E��n����}_��~ �kTΰae%%	5�&����L�׾j�V�����CB-b�}0\���9��>ϋP���:P�T�%�*,!j��tR�2#�Z�,qx�� ��i�M]�.�T�D9}�;g�(�KM�sq����]�aju|��OB�"��Z,!�"��/��F�� �F1 �X�!��ڹ �2 �y+�P���|�~�)�D�:���к^,d���.��/
W��C'�[{.�ך�A�}*;���8�dH}6��޸�%����]���?SH��8ZqL�$��?iҵ�̼O��A�R�$p�!��3��<Ք{C�t���iGk�q>��/���`�l��G����.�v�t�bAL;,��M1�L/���u#.�|t�Ykd��� h]]���Z v�+^�iD��J�R�Pr���� w�Ո���=���Y�>�=�Q�uw�`�Y��a�k�Y��>��b�4�#�@��Š���s��k����6�Qpv,�הt��M��[۾[�.�Id%���⤙��+{�=�S_���MJw�4��4HI7H��(��]�"�2t�t!�twH��5��;���[/k�Z�1s�>{?;�{��Gp�9U\�XX���M�ĤT|"�-�&��P�!��B&Uϒ�t����9eV�����P]�YDp��3B_��_-��C�DG·��Ԙ'���Y��@�ظ�cߴq���vh��J�H��ϰ���*3��.�I� �2'���*��+�����u$�����|	�uFw����Z����Y����w��D��_�^�3�3<J�|��#�yODI����0�z��������
ǽ�1=��[Jx=�������Q�^�t�!��j�*V#Z���w�ߢ�����ݡ`�)�������5�J���Dh{�77VX�M�m��փ��V��~$P" O�"� M��o`"r�c�;{k3#j+����&@G�GO����h���l��=:`�o�s���<eH}���f/8��%��`kP��7�D���7����Y��w6rE~*0/�u,����rg{�:oH���y��;�X]�\?�<�&��]g����D^�r�ouw�r"m��B�q�ɀ��Z��Aq"�:�k����[�e�LtÝ���̻�)B5T����|AC+���YHq����:24�56V����@�x�,��j������I-�~~��^+���c�?D�h��kϪ�<�x���X�ҦO�LD�Ժ��e�B0c�CR��|���7L�_8Y�&K8%�Z��A��c㙜	�
�'�Ar-`�	����<;f~9rú������?���2�@����.C��]��7/3��K���YR>�1�6=��:�[��c6]`D2�����h()b7��4� '�T~����?Z@��P���Ip���޲��<^T|�'4�x���"z(�A}�	�}T�LӴv3w�����`���2�o%�Pzg������՚���!�2�?*�=\@����~�caڛ�Wx�]���$͠�ú�S�/�f����W�\v��D�}��ێ�V� ��__�?]k�誥�l>�j�Ȝ����/�M!'��r�Eb>��W�%ф������p�-cw���R2d�I����j��^�ky�d�)��^�p_+b���BE��?r���y��$�]��.W��
Y��'�/cmiq,�;�����}��C��q5����D��t%*Y�gm@�����~է��� /4�R4q���s��a�~7j:֗ef=������k��%i'�ᵭ��8̕HZ�Pu��Ǘ���;מ����2��(�<��:t�?ls�>:�G��������hH���T�=z]�K(8�D[�c�*�i���k��H�w��g���8�-D��ރ�5\j7$Xh��fY�D�Z�Ÿǎ��/Ţr��1���a��/�ݩ��G,�q�Br���F�v�q'7�
��J�9��j U(�kz������^M�ѓ�y,H&��ꀛ#�T���8�x��S�3l�]�4���5q��0��B=u8#F��ف�i�76�ĭ�щ�)�Z/j��Q����S�Wې��;0gw>�j���8�l)M%�1h;�Ĩ���ox��kc���O^�̾��~�g>?�g�Ba\,��2��C����nj���h��}����{C�^%��:�*m�d�JI�	��[B:ʏ,�4�F3R���"�@�Tr�4q�P��x0S�.�GU�h�}A�ኌ�Xkb���]��^���{�oG��p��%?��G�D'�A�j�ה�4QZq�!Z��..�~;7W"��9������"�^�.��t�9�]�/�Z��B<���53K�	�Qxxp���Z��	�ߗTi��2���g�us�6��Gaԉ��C/����h�	H��7�T�u���Oo�m�.����I�B|���L<��_���r6D�#	�sKF��_��.^<N�|�:�sƣI���F�M���𯆣C����Up��4S��f��ܠ�����������!�;�Vaj4�<ȫJV�/Ya�o7'���?��]"'������@���P$��F���.��s����DX��4��i[.�;�G�y�Jv��@��������� ,#��2���͝/�g;{�5M��D��*�L\T�ݽ�n}���g�+�׊���/��{��~�	G*���D�ib'��Yb���=[[�/G�U^�%��Q���@�{I��ؽ�����P~���:�\����+�%�������i��eu�~��5�
8Ħ������f^����s��SW�W��w��X�%Yq��>�7?:��8ܙm�.� xߥ4�]�|w3�����?	�Exh�K��Ћ  �����B]�^W���դ��w]*	-���4 �m�����{̀N,�{����G���@�N���m����}_X����*�jSN�1��,��}�������Q�m�H��$]V3�ճ�8��<^O����tܗ`�t=>�M}��U����L�e�A�i���3��D����jU��T^�B��й�F�CQ���=|�7��ʃ���K��랺����n��_Y�]�"{�8���l�	c�P�;.b_uu��1]��&�d)��{-� �D�\�u�;�^���b�1^N)R3F>���'BHv�(��Y��s�[:���}��Æ���/����Q��\�$�hC�bo�����q��CϵAD���q���^�$�p�D��*�DX��ECL�2\�Op@�f~$W���1��I�_U�NS�ES��lW>1�~��t]��9 �s���P�{ ��Y����T�!Än�� *=Mj��+��1`0a�+%,f��]#)u
��AGAr6!�̝�`��3g��Iwa!$)��k��x���~��u���x��˔��1��� 5�s�A�^]^�e��!����f����J�����"�uW,�h�Qd�W�	@�����ҿ�n�R��x+Y��f�	?GQքJѧM��}�t})v����,�R��2/&VԱ��0�ZZ�'����G�x^�9>��c��|��¼�qvN�C[�dM���Qu�H:F�]���;�i�o��=�<��/���Y,�`b��i&ё�/q�gC�6�D��=M4����T���dm��o�I����v�>;/���%WͬX3���M\��|Ed�nLQ�;4X�ĳGGR7Ͱ��@���=YYK�{�)� ��u�`ͦ $ �kC�N���B�Њ�8f�B|�����i=ޜ���]�}q����؛��K�y�g����ZL6{�Sx��G$�2����V�:��<7п�I�+��뱐u�{��g�,n�(+A�$�R���.��L!5�?¥��rjҧ�a!':T �0��$�ͥ&��^h��6�;v������^���-�
�7��Y<��E����f`�i�:���|�y=���E��r��)�~+��xp���>�{J��_�!r��d���[��0{���d�2,�,��W��u�'�
z�u�u{�g,�B]�q������7+��V���Η0�h$AF'�\$
O�!��np5�|�M��6O�`�;��9^<CK�4s|�W(ɿ���7�N"ڽ��!�xAV"��7_�RB
8E�ذ���<�SF�TV���fl���M,�9&�{h���ŚyO�B�C�o�J�ޠ��z��?}R���1ߦ�;�٫7֌�>r�cq��$H�}�[�2�Z��۲��'Z���*:��^)$eDYA��4ee���j�V���/��������4A\E�C�$�u=��}��r�~��U�)g��,_�ρX���p��=�jsFW1�!0���<�V��s�:�0�)z����
/��*��'n[2/��o�U���pX{��D?�M�������5��Pwn����0$ M�Iy뢏�dI�ώs�;����I���Vӧj���m$s�����R�u��/j~��="���^z�X����Xk2�+nG"�a+�U���{�G��oCuzd���}-�q�	����OO)3[�%&�̇8:G�&c��~��T����
�����>�ޗĞ��6�k8�eP�\_�]�^=Ѥ��iA�.pC���r��n7�8����z-�����Vh:I��E@ ��-�i1��m^�Ԣ|W�.�D�#=����v
%��޽KZL�."YG��r�K�=g����N}���Ђq��ֵ��7bpJ��Gy��y�<7[��d�髍��Oy�?������ّʹ7�=h<�����9�n��B6#9�+��y�;�f*'�?��-��g=�cG�EX�D?{,��-�4^��lS����V��{�z�Bʌ���#�RA���0��0�?�!��{����[*F�I�2<{��}�;K�Ȓ���m��j�.��XD�5��˒m�FO��������U�8�8�".z��Mީ�ϟ�Hث�7�+��a��pn^9����N���xx5'w���@e�JE��r#���:�Xoyg�H�bb�W@V�}�Bbd������κ��2��Gl�r�>��}ƽY
��qs7O�4�Ք��y'��{���"���?�ڜ�u�_�,��Wc����x{bg����AN����>���K�-G�cq�Im�91*k3�ρ�ث_ک�e'H�	+������p�n�^�gd�uÕ�!�L�/���![w(*���g�<�S:$�����T#~��׆"�tEq�\]6����Z�&&���������� �n�����[$^��I���zK���\�[��՘H�w��55�wTz��u�@������s��<�g&'����dr��ipY��I��	������П��j�0 ��5 ^W�Oݫ��l�V=`��:B������ƨ��8X��c�L��x�⿮�i�J�S�I��/��c�g=�|�([Wf #s�:Qzj����5ir=��FVF���>p+����&q��qmZ���4��]�L/hE���y�"�B���A蘁� �S�ˬ:/pӸ����/�
sT�E����y>����o���'��}Z��tǎUmM#H*���sQ����/62�uڤ�߁��Jǳ�*2��fg=���;^ɀ%�z�4k-H1�~�EZc�Qvҙ�� {���yvf ��K���v$�/����J�_�'�U;�[Z��8����Bd�rh^��fR/Q�C?�ɽn��&ӫDC�r��^��tNW1�0�Hd�cY]rS����,c��V�>�Cv��i����j�W\9�[>c"�zFR���2�bH��k�����ɹ��}/=�O��(�zۙ����{�?9?�%�ŢgiVO.�"�vh~�\��^�oV�BM�^�5Cg�~��p�b@��&s��x��e����/�a$U�֫�$J!��oq�b��
̞�X��L�����;s O�oQ�5�R�z5�lZ�M��1��S����&lYn[9���h�O����.&�b:�f�ǯ�Bl|�);�����;g4
g�V&�Ū�" ���٢������ %>ߞ������=�yS�[JFuϾ��͸���3kf�Z�g�+u�x �����ƮT�CO���Iv��F�"���"B@KWm�gM����Te)���Ԭ�7�>�W��70T\9�����7�L�9;�Η�b�g�Gc��9��I���xv��|'���R`0�0��32 �v}�d?6��lVݧE�4�&�^��"�ҵQ�IĦ�'P�nHܟ� ��$D�(�a6U�c�O~��Fsv�����g�~��U�7#���@�?^���<��n��zw��|5�7��{[�\M駖��}�B#GiF�r˕�I��S̙6��&�ޭ麋�kS�9�ۃ�pu���I=�GG7H�+��f�+��U�0)֧�$բ?��-2:R�f�kl���}�I'�������;������	Z��r���zgv�y��;뙓�;�u���E^�(2�?q�<�1k�Ďh��c�Ѧ�	���Z��R �����Y,M9m*��/b��#2o��H_,K4�-�(��<�O拓g�`�D��!Tm��s�m��Ϳ��F��Շ�u�HV��m@�G�y�"�)2/��>�������PAc";ڻW�_G��~)�����n?D���Z�D/��������&���5�&�n�	�i;Q�M���(5�Lz/��\�|�u��m�Hg:�F�n��%�U@����4�AFL��C��z���f�F�r�/D1'h�^�P�i�t�C /"���"eq��j?U˽Ʉ)3�d�����R%�b�Yع���1��;�:����N霝ؗ��Q�������:bx_�*ߗo8R�xr�<�����|/�[}}��Ef5H1:p���~q�<-/b�!@@�gd���Rد=�Z���%܂�����J����RG�:�|c��tP��P���KX'�߲PBN�����JkQ|1�Wn�e9]]a��z�,O��@��*r�8pՕ�/k:��@�����N��jT�(�r>1�6fSI-v�����k0Oۿ6���f|k�X�:�[��^4`9�ޟ�u< �I�e��9����Z�gVF;�3>��\l�I�Q�1~��d�"��6�g���9���F�U`��u��t"��y�`�������qs!����;>9,_�כ�3����31!G�w���5�J�6-t����$xr!���*���d��.��L�n�F�x5Ɍ��a��$���فg�ź;:��u��� �M�w�i)�Ot��k/�[�a),�X<�0)�jY��_��|�k�΂]T�g���� ���=��,�_��������$W4�  ���F@yg�/��=�J�#vKJW���S�YO�-Ę������OM���]�"S��p�_J�zP��V]VF82��z.P^Q���O{��!�!1_�C������N�g�>�����]ϙ\��||�<���ꅎ_O���N>9���Y+h�l}���9T��49�F�˾g��L�-5�����e҇p��іE�Ж>�y&�ط����G<V�}��!�{]�9}]6�Vr�D=#LM�b�>ݦ�[7޾��n���m�l�	�\b�����B@��1d7;hvul��E�xܮŹ[��at�����N�� 9⯵VX�h�����&,�6�y
�k���}8Y�`��9h�L=��!Oǰ��?�%�����g^T���v� �ă� �ѳU ��Ŋm��-�����3�Q�Ga��9�$-�e�_�=G�Y�=���˧ҍ��̞��))[h�k�f�6?��s\��Y^gU�sh��ȃ�`�o����3�K���ݓ�,��n�� ]5��u�wbxnM �X��=d�����jM�x����즬��*�}�mx���2����d:���KB���B��_H�P?�#p��Q߶?��J?� �#�����6@ܾ��]`�]�O���W�ݍmΏ�����޶Ծ�?��=)c��m�G:.'���s����g\P��Pa��VrӾ�X��kԞek7�h5Ѯ�dCMw퇷�12���p�Φ��_��p���W�]'4�Y�}o]�����H�SC?�нxm���;�/p8�9�J��~�����u�n�%Һ��'1��ܚʂ%������[�P�U-�/q¡���bSدRJ��c�V���ƪ/H�D�uVCw40]^�eտyy�,��(2�H����� *1�Q���v�D����|W&K=��rL^@�ft�S��jU�뙦e���������S�E�����_�^qt�Z��0�6�Ǽ�u"^ta�d���aZ��b�+��eV�I�	�����%���E��?��x�e&�k�.̛�����it�aQ0q�b߉i���4�bX��9E@2���Yo<^�3�?@��{l��,l��%�������gn�Ռ.�	�܏Ė�����~):�#�Й,6R��Y���D�v�g��я��L�F	�آ!-�&���g\\_
�K�~��%z�h���E�Õ�/��+�˝,�}+��<��B�-��]@!{\�PuR�L:μ�������Y�xThWgX3�U97P�3�kc����K��_��WE�=���݆<�oO}}���HƁ/�n�ް�|��ߞ��̣�N��oX��/92M���77�t�/�?�4�}#�-�K����xQkaT\m������۷���1���k���͎=���{��,`����\v�X��.s������T6����w�}B�H~�����[�\��=B�� ��-������|y�\k��	.�
���x�鰐�qeڳ?�nU�u����6�'GO~�6H�����'����M�Z�ۻ)�����nة�r�����֤��n�H�y1O��*��Nͱ�#���k��_�,J>�!f��j�wn}����oN@s��7.$+��������_��=���Q����o{8b7m��w�C�AxA�|���մ�#!��2����]0�)��*��w�U�N*1���4.��H�9�+��psj����t�P�	��K���Mr�Ϻ^Z[���<~�.�����?�>�{���uQ�Ǚa1�<���>\��<�	Idt_��ޫ=R47��~������|CYA�^6{S��-r����:���B����<"K2�F��{o ��ʑu2�� �=����?#}���:�i����Չ�˯�:18s�s������S�6�s�:W��4:	Z����^���o/�iI3�� ��a7^�y�]v���x�T�[\��2�>�M:/ˠ7O
�2�#e�J��R��im�<�2���%wHg������p�6�����㇜���A�+Y7�N��cjN���͊]�A�K�L"6�����"�<�)��	8j��r[p�����NW�d��y>R�%>�9����K܂J��4d���Y5U��p%�ϣ���I���Rݬ����R��u�>������W�x���km���.M���W��Lv�"����C�8��BWͩ{Or�!z2�F���sa;��z�f�[���� ��n=r�_��PV.t��1�(����0Y�G�j��؄6�Z�]2��K�E��@�ڞRz[SB��1,* f�Z�E�<�#��n�e��"�ti�����e���,�ֱ�<�5~uws�t/�i\���xk��*��E�\�h�+4��l8h���L��qM��,1b�������Ce�#��ӹ����_�D�|�><%T4u������e���qqt���]ښ�]���ਹ�=�+=�w�&�t�������|�rH��܎�v��1���s3��m�����0Ul�����5_����D�f��YZNA�YG"����g�����M��&d
=����3B ��B�V:A׆lR�&1W���P�k%-�ZF�����C���g�+��a{���:���4Ep����+I�d��q�i8�{�5�j�XN����C��$��ꂇu *�VG��V�Y���`�\&�_W�/=$��!+(���K�r���&�X�	�����c��R���~4c�������"Vc��c*鞥��
[�j"� -T���f*Jϣ~�B��g��j�-]��~Ñ��]�,l q��Qs�0���x��#��|�PqK�H12'`�N��_�s,k���9��w,��2q�H:�=�)���Z��7dX��g��RӸ~=��<�a
���^NE�:&�^���Q9=l���r7�L�qMƧ�N��4�/��_���~�1n�(*/\qx
�d'�:�c&♡�J�<��� �ؓs���L��6�]��!��#;7��5���^���D2�S`	�k����~�Ǡ@��qջ�Oy��Q�,9�
�k�q�uO=�FN�>���w\T����z��x�$�j���_��mB�|�䇸�#	��i�(����Gk���1��aHUu��|H6�Q�P��ܜ���@�v�����2&�QBс ��$�*�7w�N2�{�*w�e�A��1%S{kw%dV{l6���%���hIձ��؋�A��ς��}�Z����ڠ"3;i��
��K�t�7����䉣�z��i{VZ'ԡChjƝm�l��C9�������gl<�%e*����N��6�ȮA���Z��wP?���A��[��1��	�<�q���ḛ��Ԝ���4 /�[�-���q����E�Si]Mt���+�e�H�cd��x��o�__rvЁ�/�/�̢w�~F��뉎p99B��v��}���Hf��Iq�v�N~��XL�@ҸG,PA�x�$��2�5�@�B�1fLj���.K��i�@�@�����;ӣ�Q���1��#{Ut B�7����7{���s�����T<���.^2�o�N�{8P�K����9����>�w�1u��R�M��M�nI�[�N�ה��?a�d�}��r��:ڧ�b�E&���Y
ZA�Ӹ����w�����Uq�~}U
�;qC��iOZ ��fN棊 �ر�~�����C�F��*#/r��['&���x��ZW�8��,������ �ν�Տ�泞T�p���Z��l�\���$@�I�X.
�K�e-c�5F���hԛ
�� f�9 �^�W��ڞ	J�A�g��Q�-r�ga� ���k���u�qS�EVРk����T�\r�$����$�11�?��)����~�C�*(����c<����P�`��Tq��B��gr\Ou��O�|��E�Xs�8O�q�B�y��5	/4�I.� xV�x���o[�Y�c�7�i�%rm~0$�`j�[�'��Iq߹v����P�ܓ1�t��#�Wߕ9��:id3�(C\c�����Y����2E��p��9"����\՝���P�pBͯ~�I��0R����Mhl�N-����������f{�Tk�i�y1�+���^^����8����B��|���L���<�x<א�Rؽ�J���oj�n�%K<L��S#\m)�ϓsH�Q���`X�28�{HLm�o�v��aw�lk]2]\kMT]A���I^��W�|��n��	��������1��f�r*�&	������Z2�tD��Rb�IN5�������d����>}�gگ{%�=�[ ���_�Z��4�&:T�^}+(�?.�$@��������_�i��B=�c~������(=Eb��!�-�<���)��i��g�b`��u��{T�E��#����]�ۖ�o�A��qcu�3V���D4��L���yQ���������m֌ ���iYYJ�=�����XJH̸�{aS���O�,Ȧ��"�Ux�7�����ѹ�s�`�5^�h���0��>�2��:&�z�|O��QFyͱ�0��豤�Lo|��1�L��>�"�ʿD�T(�u`�01g��e��T�0q 	�_�eP�&P��։v谞���ӥ'\v�:+0����� ڲ�2�s�J�r^��{��u+������O�e\q;��Q�/�pb^2�pm��`�!��l�t��"! =u)hz &���e⍴D��ג!~�R�L!�׫ut�\�,m�^�-����~߃f�\׮}�O�5��'�T'�I��cD��	�|X��NA�۷�|<�d��¶L {�M�f�"ʳ
wf�t�'ܱ̊;"��K{B�R��J��*�|r�Ǡ��muR" &�X^���u7���UIN�{R�]����J��?�n��s��
�O�m�@����qԄ�ŐY�����E�^z�Ex!`���s̑�6�T�2�hv"Y2��QBN�C�}�6��"��܄|.�H�Ӓ�b������{ۄ���\�oo�����O�5)�:��8��E��$Y�1������>!KX���欱m�5�E�aj~��ϓ��g�ea3MT��0��Ԍ /7��+B��� N/�_RL-+��YGS>����},N���_If�%�?�\#VN4����*����[)){/d{���aa�5����j���"��ɓ,"�q���g��jx��f\oSJ����!n���2���z�l&���1$��˕����\�w�\��1���d'��֝�JoJ����n��,�6�de)�yO��|h'y�08��#���N��[A9X�(�9�2�[�  ����"&��2d�g���){AX�g�ϋ}�ӊ^��+�'��.���L?_~}>�u�´3��J�8�n���i����=N�P����S���r|���ӘR����b�Z�+n�W>��l����"$nÊbS]���<喎6���-q4�H�aW�m7ܐ�g�E��Gc�DD��0/��|i�GW�:�S__^�go\�7��H�w(���+N�� ���&�ٞ�!I&Q�7�"?o"E�.E)�(��*Ðd����b d��$�	IQlQz�G=�<.OTD�2�B��t�k������X�Ġ�7U�7lj��~g��z�eځ⢩@��f���F_��}�E&�	#9���skN�Is�&t��)���M��bI�or5D�uJdcɔ��������vf�c蛼����J�?q�Tr���;D�q�"0�M# M�
ctLX�{�7r��PP���.�s7u"���h/ַ���"���ζ��|���������#��\�q��]N����#���`�h��$\~��wy���h�,z��K��+�����������R]������i��[*��e�����m����t5:&�pºl�	S�wߺ�a�U'�u��;���tb��w"��o�0�e�8�F4S�UdQܧ�y.�j�5�v�m���"[��.{@`ЌYg"�r㵡��z,*�l)��(]ٴ[Z�c{|k(WC�."Ӥ�x�N�Pܔ��`d21�u�_|eśG�K	����O+�#����\�eR$@�Gz>�k`hEI�e�S�D �Ҟ��4ʏ��A�ֽz�j�I?��id4.1c�ϩ�!��`'�ۈ;&��٪^������b����9�F�7����?oUL8ӿ��:����'��ʐ���{����B�%gS�t�-X~] ;֓(;����m�b��V����?>L��F�h�bN�ޟ"�;�D���!(��GLB���wh����6��S�6��=��'a<��;�J�n�qn���l���oٽ�gYrڬ����+s�7Η0p]X�^DK�b�OYB��L��hbyVxw��jU�W m���B�r��N�������.�5�*h7���p�Ԍ��̦��_��!�W7���D�%F���<��8H�Ř^��wd����$�F���gP�wC@_��>���>���+���g�z�a,?8�fn�C4���T��ɌQ�&��`�_k�N�caFZc���`��5H��d�C�dP7�t0��l��zRR�(IMȠ���bԒe<�}��e�x����y�)��k@�Cc� ebT�[(�-���Q����1�߸�s�_f��F�lmkL+$��
!I�U$�%?���9n��E�\~E���������u�{�
I
��}I��A#����@i���8.83��\%VP�;��(�[�=-��}ǥ������g%�C~�CP �ə��W_ߘ:���1�M;B�"��浲�������З���K);Ȝ �I�c�UR|1b������y)-�|6�#ʠ�����+Ln��u��z�M�<]78�"� c�;n����<{�fU�����iC�l�O�+9��A�2J����[���U澂2YD��٫��!��΂��({�8�Wf�
��In��L.wk������Qz�l�\�%���1���p�����{V��q�����0�AS�J����:=-��vo^�掐���J/�9
zƭ�5 Q��1��!"S���$��X���-����@z���ixu��y@�xF��HQ��f�9���i�����u��1��`J��ᩇr�O/�Kf�n��Hi{n�C�VQoA���{4���&{;�I��F�g�Q�- ��r=y�g��Ss�Xw�$z ���3���U���e9]bQP�i.�F"��X_���
F�\.@!t!#1��
�Hn=��T�&����z'v��u�����l?1u`�ġ'B��r���?��r7N�ag�DYy
!�XQP�� S�=��m�x������M�=;ǯ*n�A�O_�_?I�!9�T@I0��p�o+�(��VFp�KV|����f}p;�V)���U��饧�N��ۣ�Җ}�[�@��[~�K
mB��Dom��1�����pX��8�����ܩ]wgu�g0��y�1���¿r�=,욓7I�=��MҾ�@��E��Qb1p�߹yx�W?��d��&�7��m	�L6���|C���a���g9�������yJV[���$@u���M����
�M���@]R��q��rkg/�.�dKD�f�"�9{#蜢4Yad���x������V����M�L�X�i�����j�	O��f���4�����bq&��D>��0o,��;�O�� �j�ܘY�\�a�'��A�t��Z���3�}�wP��Rq^�i{P�P,��p0���F�}���vX�X��(����RS��չ��S�(,�9�������� g[�e��V������@S�h���ow��G�>���2f7_��>�X�;�$��t6�П-���=8��X�G/qf>��4L�l�|wB��#��ړƹ��e~�L�eC'�w�-,�M�?L�}�h׾;f��0���F�)�f��$�k�p�F���(���\����?�{q5j��k��턲T��$f`�P#���y�j���|��#� �*��4�������{���{��ʿ�'���U_񽏘ߤ?As;cۂ܍�=�"��|
j���|''�шZ�`�?��]m�m��Ȁl��vc�$l��8}�K���ٳW�/�<.�;�ڳ���W����U`� ;�����P�ُt��?�E�UJ��xY�V��	�{`Tb)��}*x�x��~:u���;GĨu���y�������U�O��Щ�P��.+Sjl���75 3z�D)]�ҀN߶�+O���2�T��b/s29V�W�T�9	�,�����4T������kF^\_��X�4���--=�S�b�����'6%>1�ք��|7�d&�L�$g��U2[�j ��P�����,��/SZ��"T������h�o�����YE��H��OJ�'y��'����}�=՛I>�z쩔щ�L
�Z��-�ў���`=|T�����vi�s7�*ݧ6,XCn�L�t��>��MO"������M�@�^�N���W�������@��3�>sђ�l�a]��:o"�>~����;���$�v�6	3����>؊�&g��=[�� �B@��Z�����3���}�,L���ѴM��D�K7��N�$Ҫ�����^3���g��t�a���-jӐU:SA�T�V9�p���
-|�,d���"#���jA
<���\��aGc��r�vW����2#�԰m�4v���{�o�9�3�L�􉐆���h'+XM��3F�'�|M9JQ
�6�07�������uyjƦ�7qO��;���6�,x�w���h7�S������}�>5��7�*[/�i[ �c��buq���38�[v	e��V�B�J��z���-��[Nh��2�]s}����6����CV�[����HA�t������ڕ�t*��ܽ��3rp��Vh5pX�Uޣ]
�"����q�a���'/����Dj`,җ6�>B��+�^p�ZCX��:�/Hi+,{�� G����n^_�]gbr�!���k{KPv�I� J��r��b�\�v(�N����_�~��=��:�� n��~�2>cם�����2.��=�9�%Tt��g��IH*�]��w��� \7Zwfޔ!���ܠ`��,�W�f��;�%���ƿ+��@�����S�b����]R�T&j������~5���?�l׎����Q'5qՐ(+ث��.���� ��.SR�h�=�v�J�ր��q$���Pa�z�=S�Q�>�O����]_���%D��3���p�6�w˄�y�O�v_ӮvQt��&���x%�qڧ��;��D��B����1^<���g��]WQ�o"�n�s'4�,��f�gʢ����C��g���׊i�)r���G"z�h҂�a�����9��l7��"�a�B�·����D<l>-�ZO�x�Ot��V��&},�(�s�̦�{�l���1�����)�HE5dp�^��y�N/���k�g�wyA�7N*OOe�<����Y��r��r}��_sQ��
��C
�C�.��ӋD:C�r�������|Tk����(	�:��r��UP�V����pY8:���3�����8g�ٽNH��5�ۼ�|��L#�dQa��&���{(��<^�f��]'�a%!]y���ϰ���	������-�S�w�����a9\���6��>x�	�����0~��E�{��*��0z�=Ì������̓�i��b��D.'/\آՖ�+���S��Ŏ�b�E�J[�~�O����&�wT�>���cR��,�8U��F'��3��op|X�����ZjP�u�>lVK�W��ꚹ,�&��Q��ͧ�NHv�[z,;m�Id�eao������&�a�p�Ĝ�LXn~^oKѫ,)W���!�_B�>x��Pݓ~^ +/̩�2�!~'�xu�|8�6f��ʎ�"/��	�Y����6��QU�S�WVF4�82?���԰�\ۀ�KM[ぶ7��>��t��g߁o9Y6�h˦rpj�B�8�iWE��� ��Rҥ��)!����݈4���Hw�!�A:!� �xo��{��χ�f��{�u��5�d��)�`<��������m�ý��q�3���J�Uk3͠��9�z��{joJ�C����ҵ��˜�y�=i9��,}���5�'��nWm1��\Ȓ F��tq�!)m�ǣ�(>�}���d�^~���_�1��4�����侸UfYb��s�t��ࡐl� ���iڕƏ[���qI�/f���U����^�����9����^%��j~�5�z���-��ⅆ�&�
Շ�˶8J��4�b2��ə�'3�6b�'�hB�H�*�ܳ
^Ֆ�6���ri�o_�'���V/|^���:-Ȍͩ�� ��XC&��қi�sd�V~�e!���tse! s�FI�}E_�K/`��x���{.��>����@�a?�{�a�wmo)3�p��U� ��Xk�����q�Q��O���e�	)7w������s�A�@*�}*T^�gn�X�R�V�zx����X>nJ���hb����iÌ9>��R�3pa!6$�/Kl���������v�]�!ۏk��x�fb�t��o5	�}n�e��%�{u<�DI�E.���Z?x��~�u\���v�Y��H��w:�����%���$w8@1�\7��xO�#�l������g��*���sx�SV|���O�����)G�z~�v%��=����w�M�+4��Ѹ�y�󸪖LN[)���_A/���IKO��rs���[���&�p64z�m�\5��A��M�� ��[���}k��CEw⭷�ɉ �/w�w�z-SdvBض��8Ɯy�����$ǯ��m�d	�80##�P�5�;�![��ȍ�I�����{�C�5�V|N�z��qZ���v�=�Z]6=8�3�DN(*��P�m��YP��ТI�$`<P����E+ɕɶxDs���/D+Z�s�E�i�DAE�R!E4,�u��x#��q�F�P�/�"m��# ���♫��^_K��6��u�޳��]��4����t��\J�f�@���Jy�=��!�0NRw����ֵ$Y��_�SLb�X�4}�U�F�5�C��4� ��H�h�S�K����2"�����̻!��bJMA�W�DR�X].ɥ��}~��G����udF�tJ�3�����o��ʂ�[g�M�l�r(jH��u�{���R��[�A�q����tK���Zq���L��"���^r|HNeR`n)i9���^[�rF8~�W3F���O@3��ϣz>�&���h�J�k�����{ڷ�7nc�^��S/�?� �1M�p/�+W:Vet�r�)�\�_����@]� �.HW��f
� Ɲ�4�h"&�JFP���X'�n�N.P��h��g�Q�)�0!��nX|��$� ����Y�yc��/ЙַK�I���u���7���d�����nQ@�]d��~A1,'�̓�[�6�*�)7�r84�<J'O��i�zw[|�-�T���'��։Z7����0}��3j��lzhY�:��d1ׁ�����H�)�~��YPJч����5��;E�?ۃ��g�CG��d+W�#�Z�j�ܭ�Xl�_�Y�(h����`lC$:=���lG���o�}r���O�`�%Sk�Sw���~�Iq����G}R���5U������7kR�i4�q>�g����2�Kk�I ɴ�-ݸ���,	3n ��t�+�1 )HU`��]�EV�#C���>�<�w����hl�.O\��h��̭���5��낦K?��n�Cz��v�F+�c�|�%l3�j!M��`m}�����rh{�	q������9��_��m�t�o��IB�{�h.Sgu���"c�����:9(y��C����ADco����Fd�?��EU�j��e�TS?���\�3��⊐>j���[�ނk%��J<Թ�]�6<���<��^���#�� ��Ô��~ߓʠ�*��j�$U�w�Iʥ����ir�CJ���g�h�+��b�ݣ������$�N�rV�c"jm1����8~�Q���I.|k\v��^8�����[+z����f�+x���!;2�PX#��~B�1V��P;"]~�ዦ��>;8G���L�wAq�*�)�
WU$3��ϐ�Mn_���Ck\�X�-���}'ᑆf�{������X~��E
�Oƥb)�K��(~d��P�����S�Ū�.56�\��/<�T��8�]��>����T�a\�5>�2����x*Χ#����91�97_���	ڒZ�����)0��M�+[�+eY��Lб9��d�����s?:���km�w�IY*�,����۞:�o����kk�+s(�8|��,m���]M`�ԉ����<0g�)o&�sm1�7�J�"K�S���!�6����E)���� �I�Ak`�1n�࠯�؈�_��	�3?�7)<џg2g�Q�]�����SHe֟��)U�>�f�(R�2��1ܷ
maLvűkdr��sy7k|�����ʇ�%��XN�R��!H��*��5�,��x_L<y�?÷h��-��4���D'#7$/��U '�_h��~�7�R��݁/�	������`���H[�j��b�	XZ4��<��%Ng����rA�=`�WEqt�֩H�)§�������d�uث�_�9h��!y����zq�zICC*[� �jgU�պ�n��&R�^ ��6S�o��e�є�;bg�S��x�L�?S��{G*��M�����D1��ڇ2���m��熪�ǩ�4B`�T��=/���K7�'���	�,���4b�kB�D-8��&>Ӯ��	z,r̄C�M�F��-eg�Ζ�ҧH"匦T>$&��ԅ�wSb:��Yh�)A����/�DU�,�u��SL����J�΋�=LYT��߂ZN�Zf���R$�&;��@3���*�Vt�Ow�cSV�=���*��ݳ�����붠J���	z���L�0�IF�\DR6�P��N&@,ж����p��|镥Q��c|�71��|�Z�'1�X�]v��HZ�>Py\܀��_/��a�a}lK)�v����G��h�:��ƄQ�4��ԧ������a�:wMJ�O�
���\����f�0�����\[��������v�A⩔}��|@�O>5��n�w9
��_{5����?F���k^���3���V,��sX-�h4#��d]O>�ի�m�~�Un�w�>����tTK���l;���D����'?6Dѯ
�h��@j�F4��x �*b�c���:�
E������P��	L!.��[K��`��%�a>>���>��aSX��t~�PB1��z��ka]A��Ok��A���\��6��N|ѵ�{�����8��$Q������Y �ΰ�39E����o��/W�#��
a�cE��x�b�s��X�ν�S��*mWoa��jg^rC�ئ#1qL%D�V?����U��n�^�W�S{A��C���;�-���|#+W�b����^�=�U��Xs��ۚ��4��J�`棧�N$���Q�fh��^oxBZ���l�ȼ�V�ү�*�����MN�#�a��ǀH~��>�y֮�'D����`����$5��q���h���X��+�_#H�?�z��M���a���sO�(m�$�&�sD���FtMr;��Z���N |�n'�&���yk��fCFA�E�篝�%��|E}�׿����e?���1P�3�<�K�f��k9h�!�kZ*�5G��t5Js&���z��_L�YY��4��ǐ�kME��kɗ��=,w�F7 ��͜]�b>z�����CNN�Dr��UP�9�X՝SD9	��wz���Z����Vw��,GAs����,F�SHNB�C4QGz&m�Te#�r��虥�jb�\�*m;֨M ����[�2�f�D�{�/�� :ֿN�wS����չt��O\]|��:��M��.�A6ҩ/,�p '�8�0H��g�ab7
�<�J"9�R�^��iF(�d��}�~$˔"p�	9=���,�r%��]��cc�?�<󜽄�ۄh������#C9�#�Vx��ި����[|{#��&/P�e���eΧS��^DK%xфP\�=��脰y�Chrۓֺ�����S��}HX]6��g��﵇f�C>F��#Oݱ�>�oH�6!H����v~wON![yQ-�%ͭ�"��G��|M�uBqyvp�up�p�up��q�Iqy�p��qxH���eE>�B�2Uԟl$n�a��Į� � //�+_�>Gn᠁�K	���}�2u2�Jz��X�2_��o����}�È�n�v�$�gz���S����+����t�#��,,�{���t���D�	�������ʷ����wH4�N3��5�2��{��c��U�����l�o�7498B�#���7T��D����ߤ'�8���?�(�[���D��nHD|_��S�~}*�c���#��d�LqYY��f�D���Qqq���OA�,�Y�X�XG�L���IUg9�6\\\,��I84<��}h����'bbF��y���!}���v ��G8^���׍GS;956��&&�Se%�����U+�Q�Ɔ	�,��S��� !
,	9u���i�͡��u�����ke)b1a���uD>������d��4S����/*JJPs�H��tӸ=�ub���,�À0_�qN4{�ѡ8���L��0""���i�0�!!!������F3�(Z+������do�B(2[e��;�(H�go����j4�"T�����F> �1��Jyx� �QWW��A# "�L��.������G߻�ߦӳ���V�a��^�03`�x�u�c�<�jf	��M[wmYsLJOGNFlZ�)�j;�g��g��n���K�NOO���C��R����_JF�?�2qr�)(�Ƽ{w.����MV돥��j�S[6����M����� ����א+���6r0�̾y>��ݹ�˦/y��=/�������lD�lD�+{�L=�\��L���WWWKK� ������
̊��hق�[�?o@B����1C���{�����H���S���	�~�ͭ�d����D���?����@���>:�����l���Jjk���݋L��fd� ̎p{��(|n ]��Va<:>>=��(r�Nkggw.���a��h@�f�{(�%���
�tD���F-aC)9�TOSP���������P��@u@@��o�ί_�p+}}r_?���瀃��ϥުz����i<�?N���!@ )���:y$�:Y��{����N�Xԍ%�g	ǩ��2
8f���y'q'	ӻ���x��?~��$H�W7�
{
AZ��pʖP��ǟn�~�������}C-�(Q���gسN���`�?������͵����!&ޟ�P��,\�x��7ر���h������*�������?[�R���:	B0���@�Bֲ`�
�V�����|ɘȦ�'��v_4�PQ�sKw��O��	�oC�*y�����R%���W��V�dÅQ�����OQ������/������1�cQ�o�\��c�����ƋKK�O��������7k����������	���Dм�ڳ�����L.�yް����@� �n���Ω��da��nx�+�����mGqv'4�0�ya3r,lH(}ښ�։/uőI�����D�c3���ve����O����=����YY�jb��o�S�������#�jo+���b�LSUؖ5�k�Ix�"���EK�V�v�E���|Bq���1*ro�k5C7]�=���{*m�x��@�oOw{Pك��8��U����;ǅ��ʃ�|zv�Bl�s�	B�^�@Z����ߌ�\��������z~2��� �}�
�.��m�}t�AȷVM5)����JN�ͣT����A��88W	\eD�l׭��QNZ;�3/o;Q9����ĮT����hVd�Ƚ�&�([)����O�.4MŚ*��v�Յ����5?ݎf3
?���v4�������}I��H5�3�������L1��_���a��Z"�� ��AQ��W.zy�Eʕ+@��8*�a�:��}�S���'+:Qk��8�B��2�d'�v���\7����4������[-z�%��Q��x9��z S-��U��J�jҠ%q6����j#7�����w��B��NO��4����wI\پOٶ��n�k2]ukV���ϭ��8`J[�p�y|%ߓ��a[�����6��g�b��UkF;���-z�+�W%�G��u����'19;�2��r/���@)�~Fp����_��C? Q�ld�
����)�BB	������X�˒J�1�5�h��r��3��K�`h�X��ٓ��뱕[�l.���0J�5ۏ
�|�M���b��WpŊH�g�>����z�Wl��W�c����\�H�UQ��Ǆ��﫣AWH$���/e|���O�2�N�����y^�=�k�s:��-���-\�W�.�R��sO��	���C�oa��m��Y�yģ�I����ȃL�O�d�*���Lr�C��w{�X�G���e�e_�f��^?�oU�S��8uf��_��A�*�g�$�G�=�Y�WW�(�b��_Q���b������]K�������5�����b"x�.��]��ֹ�L�'i�����%Hh�}���{?A�� �<�U�U� ��C�����m��$Yb�bq��.UQ�-���oj��\��m�;S��ۋ;c
1��Ggc�����ݢ�@�YX�O�;k�0�8o�{��j�%��b�;�	&?�������hێׯfr���ؖd�V��7C��AJ���ˣV*2��n��OJ̾�O����t�\�Ο��FJf���-&������s��Ժ�/#(�E8�;��N)#]vA��V��7j��bb���9[���̄o�	�/D)�nQ����/GF���&�b�+�p|_ufB!�����/��{jP����F�N��M�=��@
�JԵbi�<Tx8z��Ik$�LٌQތ-�W���I�O�.h�S:#s�VBt�*�Ga/و�)+so��G9������K�K�N�j�{�ߎ!1�6�$)o��B��&n�	�8��S2�ˬs,�;��,X�ɨ�9�{��.-�:݉�:KJ���|SO�y�oR#����w��k����x�i6�C�'̂��w�^�a�!�"v��G�L�ρAa��J�r�u�B!����m~۞�c��Qp�_,�E���Ͻ�T�ׇ��~��C�%��!�*�0/l	m=`o�L1���O����9���>U!���{�83r*�F��a��ª�1H�6�(���a��
��o�-����HT;�o1�v�]UJ5����~� L��?b ho]|{�D������ǭ�1k��"��>)5=�GR&/l�A���`m��P($��>���V�&CO�,1X����QJ
��ŴCd��k�\� ��I�EϹ|/v�r]�du5���uv����&䱒���pŒEArW�w��7�]uH��lël,�p��ת?�����иO��*�s4�a�S�	b-�߽Vlקd[�/+���듧�MND�rS��U���q�}~+����i6��Y��I���5邥�IX�4S�QAe�=Ŷ���U��@V���FDe�az��4��M��^�����/ì4#ף��IxY�7:Fi�.�1�є����
�7͚�$z���\�~�~��i�"|��j#��^!J��{V�<�>�z[dB­���l��m���i�0�,%F������f1d\4�"L���*ɳ�o�>�)�?h�ɉ�}=J�7��?��n����f���FC�f<϶��R��QNi�ӿ�P��Mv�9�:��f��;O��b���u�s���������������<O�T6��}�����+r��yn��oIDmi�bX����U@%��BڜB���Io3~b��TⱈM�UB�㶠�� ���zrq�5�̋�AJ.+��i�F�m���hx�)���ZXH�x��F��qAdȪ��Aӗ{�1��8{KǷ��*{��ᡢ�:0n���>�~�g75]�
R�"�H�����V��ʐԙԘQ��}�Dn���cE�E(;�Xo�&utO8�cC����g�pfW?�g��kT}ڋ���e�������vzT�~� "NF�-�;��:[���s8�}i7�2p��6�r�0�&r��Jo���9Y�ժ䜃6�V;���e��ɺ �?���ɰ���d�f{_t�\��v֏���]��B�o��	�aD��7�<64�^5/U���/AT����Q>��4�n�Q����so���{�۽�Y��yM�A�G�|

ٍQZ�9�p����+�������r�0�kĴ���k�����UZ2S��c�i�z�wuՖ��;Ǘ� �K�5DsgmZ������V��Z�1�Lg��q�§�Y=�ݵ���7�b�,�V�˶�6���
�5h2
��HȜ��`���m&�����¯:MWR��X���z[#��/u��>�F7�*b��L%*�Y��ȗ��K�Q;�3̹����c�]ow�mX��3=*�q���4��8�Z��Br��_������2B���	K*y��W���tH�vn�p�����lm�=-�t$�A�B��gF$��G-��)�˔M`�%�J�K��`�a���}Q�O_�;���`�/f�������X}9�&4��EP-�C^�T���d�]#�k�I9�y"�ft�k�ר	v�27�v�V�Vj��^��gaۖV��
���;��fM��k�Y�,ms-��;�GIԇҩ���_o��b��r"L�}UjX��?B�/MueԫMF%ۯ��V�sn!�w1���l���ĻC�X
���A�Zz?��r��J0ju.���}[$A�[��חV~t+��:��c�?��,aI~���N4Ϡ�� ���mB�v����	�&�)n�P:`zo� W�.��f�ȟ����C��=O�#%��sD������>.+h��R��(-5=�vろF���~��Z�N�����V�zx�K�]͛C�;
�M,��sn�U�}(e�i��]�;�}|���Qn�������{,���� Ij�!O~��3��v%ho���P�N(�1��lh��'wI�O(�?>TTE�m\�u�����n��⭫=ap�Hox�8��y�����oT�g�ˠ;b�w<n�q�=F�q��P�����&�:�;q��sU�;b��Z6c�ύ�OL�SG�}1�n�>M��=ȗTՈ�'�-y2#�w����ę�# Z��m0@�ӓ�6B-Æ]�D��gk���s =`&���x�u��K�����s�5��Q%�P�\�w1g�v�}�5H}���f��~� I����XU�|���l���wa�,�ka3������ۃ�	�J��C��ʮ,/���b���$'��ؕ�Ƴ���Q>��*�?��B-DL�����b�jͦ�H�)A��W=�/!�����|���H�=����F�ط<Uܳ$A�:8f��xWd<~�R;|�Y�6e5vy#�&c�� 2>"P�T9<�dus��~�s,,�HS���	���6��]$H��~��%j#�\{*]��2�}�������`�3�]���v5�f]̚�x��ڵ��\��跒���"OG�L�on�=t��Ơ�_ZJ�r1��XM�s�'4�N!�)��k��"T�MOt�ٕ7���
E��D�g��ť�O��ku��~�����0IqYu\6�\C�W`�69���6�k`����(���6�x�>�gћg���ލ�_�GFd���I�꩛���v.Ծ��xK�vUs�Z_�쩋�'^OL������'G2u Z"}^K����d�񽤛B��DTan{�C[����sɡ0U��wX˘H�w��Q��\	���#EV�2�j��d�}��7��;�_jti}���@Ŋ���l�>�z3�#@�#s\�5�4��@�?V��Q~Mh�/��`'��ۻo�!c�UQ_��K�x��dV��
u4Hs�|����S >$_ ����aYi�i1�+��P�{�Щϼ�E_۰N��T���l�]W��K�����|����h��������/j�v� U/ ^��嗀_���}(�v�|��;`
����t����(�v�<�r(f(�;�3&�,k��X�{J/v�����~|�!��G�9�-@���|1=6%�F�z=f0%�?(C�!u[3�+����+�Y��rH�>v�HB* b�����Z��`��w�]`�M�6^fKи����x�e��d\�?j;����
�F�����|���w�41^u�
��!4bi���q�n�e3	/`���.p����(�ȅ���)��5���Cwr��JS�y͓�� ��R�M[�쮠W�9�g��]��Vވ[?�_����&��-$u�g[��&Y+�����d���pm���"U-v��;�s�W�G��u�p����y�3%F��5Ty���o�Wh�WH�mcߦ�D�(_�4`P�¦u{��	�B��	t�I�8�LN����PQ��oJ*�zG�EX�yP~d�Xz�E��6 7�|}K_<i��Ms_ �Mɢ�G��ԝxH��|�,�~�{T{8��)���H���)�s:=�nܞ���YÄ��"J}�����#�_��-�{��ag�l}�Mz���c��'��$�3H� ��˾�����t/RNl`��j.�	��RzHo�V��TY�ɛ�8s��L|d`�&���#y(��.��Rf� Gֽ_l�m����P)!-��#��9̫.�b@+��st��E>�ggK8y�NPnpK�Bd�a�u�����N��3g�υ�7U�>�v5&�~=GL܏�tڮ_��Z�,�/7�2ҿ�.fU�� *���vH}/ME��X���C)BހۤjaE�� �Y6�&#�yMW��S���S�9>)W�s��r�#�p)	�T�R�����n.�+�����HKg�o?��5 �z��2=0t�i���Is�%��gTb�<���W�p)�j'q�����q�S2X?G�+��9#I���u	�&���6�K!���g���!������Tq�=�Xl2?�dd0l�z8|�a�9�b�~6�fQ\Ŏ��T���7���4�q���n����Q&�Q���'�b�ۓC�i�Nոɲbh�-�L��z�ޱ�U0��q��A�H>������*(ᛠ-[QN��Y��z:��k�%ނ�[��GE�����4��1텘?�8%�-�\��.�d��p5���-2��"L����h�텗���z��5|_K{��g�ev,`�]#� ��%w�f����L=m�(��F�Ȑ��7�V,L/����p��Vt$i���/;kis��;��"f���O�����0���m��
>ݩ��Qr���8�j�+�Ҏ�!*'��)4�=L(Y S��XEq�5mV�tX,�
.�+����*L(�\�͔Gr���ᒔ�&�~�M��j߬��O=����A��wv�d����֊��*/6��bUƪ��+��<ai�FUK��m��x��T��g��s`�B�ް��
;]`���H��ݶ4&��W�(u��Yo�U�Jo��|Q��4*kx,��:Pc��l4���`1�CID-�ӥ�{/s��z �ec��$��^�������~7N��>[I�!F�O��G��n�	w�[����j7�����\JF�Z��Q~���i�����zS�EE�{�F>9�ş�)|޿�_^�����1b�eڻ������Yz	NG�,87���ѝU�0�,Q��!�xGm��5�.5�{f��لɅ<f/b��M��e�L�#�|:����H���mZFb~��̔|��U�\_�U�c�}���xl�h�@?�s�9�w�G�d-yX�n�iim�2�$�z H�Vc( ԁ��Udͩ�K����C�3�i�ݖXK�}8���|�:�Ƀ���)W�̽Dv^�L&g�*VԈw���|�������ց?�ht�گA2�ӯ�t���}Ld�Ƞ�e(��,��\�03�o5x��o��
m�N'`�~8s*9���
��O9�3�%Y r���P�Һ���G��!������j+# �>JC~6-.��D~�(N9�:Y]����q%�.�k��<��t$�a��I;=�,�"�Iz:���62�_/ME�ΠXQ��hse���Ҩ�6X���)���q��*�l.^��:�n/{��:t�l{X�V��~���AX:�;��(�R���b��b*@,������H㕪�5�B��q�����]α�?-euܖ���Zi{ǩZ�P<Ӫ:�<�A�����rܐ���<�&q;��6���ah�$�-�L��.��|xtM�� q��l��~{�h�Ёu����;��%�垑%[�A��y��������,���âMJ�^ّ�]A�Hyn8�U��VJ��V��@{V�!��k�Uw���3)����DA����{�L�#��Cڀ -��SIZa�*�`c���΢��wT~|V#e��M}n?�	�n�=fT���x��&���[c�����{��6`
�K	y-ᅎ[�dh�N���lG�}�l���Tbb�T��9��z�I�S�Q�^����S>W �S5�׹�P
�J�ϷҮk5��jY��f_O�v�4U�\�R�@��D����p^���V��@�N�$m�P]�V�=4��d7r(4�0����B���~.u.�o������qe�_�YU�,�G��-4��u���vӮ��*sT �h��N��<D4���4w`�2�9=�=[[o�yGkޛ=�����lE���)��Y�8���`�Y�ї<=��q�R�e���oo����[��� �u�����5����[P�	�}.۫3a �U^X(���I>���>��J�[w�w��A�)��/'(x'��GV�uP�q��"�t�{+:
��ݟ#N��덟Y��8-��.�xX�쫘`E�́�T}��.2��$y~w���g��_����4]�f����3�ly�"A�B��G�_ZÛ*Ha�������\�;��zό�8��snӱ<��w�ok9�Ϫ�.3ԩf���s6U�0�(n!U};|�}0�'�����?%˗�>�z^�/}���_�~*�I}�'���!)p�L#P��v�Q̫5o��,@F�L�4�kT����wL~����fD�1�կg�n��֟����$譽�G̏���(�!9��4'��o8��h�t[g�_��4���A;���̬7�q��KݔE|{��r�ekf~���w�d�>�Ů�*���Ա?��IynO	��rr\�\��>����p+b�:X���$?�#!�o��'mZK�;6�ݬ��>�	��AAP�3bo�X_@G�-�[Z�#0�	
;�a�<23�}�uֵ����e,�!��mv}ݷT�SM12�t��;�@>s$t��U���W��Q�!J�_N1#`�Іs؄jM �&.?������P��y�$ӴM�T呐�f�bz�XMT'<,�)���spqy�iL�������Z���\��F�Kt�<9I��r���py@>=( �<���C(B�B-f�#�?�O����d=�0SC�Aw��.n|O�/��^��x�_��<��)y�N����߁4�ͷ �e^��K)M���$��>ى[t-O�x�u��\)u3r�(��EG0/w>\Kߦ���E	D�g�{�gl����v�����˞�Y�ϯ�QH���@���;�dN%coߗeB�n=&+��'2OP~����!u�u8��5��h�bO> d�7Dɯb@�I����RrP�\Y �O܏�8��-��)hF �ah�f�Q,4���/� y<�p��4��;�t�=i)�J�&a�c�Iص9X�;>erт�ψ�r�+jdVW;�3��k��̃��c��֓�$}������C5B�ɣX��U�Zc�;n!쭐0l'���pf�4��\�����m)DW��_��ŝF��IVV��\�ޗ�1�V�V6&��+�ʦ��ё����M}�x�ή���s	��Cߧ[?N=z���|ʝ���R�=R��k��Z��'�lj�Wo���B�,2Z�������gAF"z]	O�M|#��bb��Nѡ�w��T���tB�Ne@7���y�y�J����_����%�y�$�A�F���r��J�NY���k��	��y��(�|�޹��05։�.l�-+���d(u3��y�����]�X&��5��R��3	�,+m�.�^��\�(E�$�ᏃiP&�G?�c.GeU^� .���,�oeW�?�XE'[��>�"<�$]��lFu�5!V�����3s��Q�T�3��&w}��XqA�
�5��(���O�p���/D�C޿�{��H@g�U��*ku3U�)�p�{!`�tuE�ཪ�B��7��4epi����֕RO��R67�9� F	D��Ng�_إ�M�w��)�s> ��l�l�lU~�{Ttr�9���O?a>��i4��w޹�����ox{�6�ILH)���Ϝ���N�X0mH��ܵl:Ơ��A�՝��"'�Cv��uJew�	oe{�+8Գͨ�W/ڐ!i4Ee+w
i�lKE,tZ�X3�b.��d~;?�E��+�iՀ�n���г�.c���7���%���DΕ܊�[��� T�bC��ۛst{)�Σ-�ɣ��bVͻv@���=T;]�P3���,F�~���D��zKj@(�(a[*�}枑��4��u�6�ڨ���q��[�[<UU}�W��Uk0.��db_���
�r���.�,Y�V�{�\	N�m�<3�B�٩�uE�f�]u�E�Ձ�m)-��j^��j��rz�2X���f)�徆�J�BS��Y�!ȥ��5��:�evY������o�C�G�~N/` *��K������b鲂|���?}��� ��Ș��0���]L��n�,���ti8ky�����#��-��L��ڂ7�vmq�5�3`%����t�h�QB��bcc��Qe�a!�o`�GT�+�B�����w5J7ܟ�hn�?U�j�!��_n�!*QmG!��M������g���>�v���E�dx^��!<�h�U���e9�sW~8f�g���s����z���wԨ��w�����s�w �P};����J��?��+ ����r"P����B���=v���󗲡Wc�g�{�o�����뜶0�������@O.�����L�^z��'��8�z`*�S�����({x=S� ��n���A�8�<��Q�j���s�'����4,�t��9����B=�f\>�A��jW�����}��l=E�ͅ�J� �BtW�G >�ӆ� 3)��ad,�>�<�����;c�UvDw\P�C֬�v���#��l�jbU����	�֛�H�3��������ʐ|�a�4�]ӨZ"�Sǫ�ܡB������	v�����gbk�f�<�l=�U�����o�B����:`1un� uR�k���&R�	S7�'�D}l(���Z=m����E[��Ө��׶�BO˹�UAj{d�
Q�)��+ӭR�����(۷J�o*m��\y��+����J�$z�c4��s�����q-�V�/15+zI�%{�`�KY�&w��h�!�c��^>F�]iSR���"1ޝ$߂3����۝ԟW�J}n'H���Y�'��4����%���K��FDsT_��v�(�-Zd:U ($���9|S�X�`���u)y3��Ӌ.՛.�ԛ2A��?�T�-�Z�#��1��ݔ���G =a���>��;��jՏ�����B,e+vբ4�r;i�@ �[;�Dqԉ�hZ���y�����\�g����_��E��Y}�ܧLy�A����Ν��	���r�SZM�8i�!�M�+�{ 7W��zH�����dm%}��lO��4��!x��l�(KjpFx&��:��7�>���{���1�v�����tM��l���_�W>�l�Z�+������UE3��+�z^�����e�䳀Z�����'���S5+�c�]DI>�Z�^X&��*;����>*2�D,��#,@�G���b�K�^�3R�jn���+�����Р7�4����[�o\�9�=���7��a�l�eu>�rGu@��8�k���a
f�f�=��:��̗�,�5O�D��sG�22	��;���N̿��Q�I<�q����cS�]��! C�[�&^�f21 ��}��J��Yx���iC���=ĖBRE~�>(B>.S'54��;7�ҹ>�ޡݎLF�=;3Q|��{H�>i��B�{4�	w�X�c���|�/ff�Ӿ��RZ��n�c�_v�����{�;[k�AU����� �Er�}����¾�ݮ�|QvD�{����M&������1�M��� �|��j��Z�JX�ʗ`c�K�H�0�i�ќ�sԌ����W06��&�V���G��`����F���:�'�'���0�EA�*��ƕRqv�%��DUT0#�-H����/pE:��E �GV
X���5���O��t��ֿ%�����U���=�K/8xz���5Ptю]�;�r���`T�� A��-���ޡ�W�C� �U��k&�'�p�Б���(��u��q/�ˌ�+�Bژ	��Z����gx�4����:�+�`*�j1Z�VXw8u#5�n��ϾO��
��ϸ���?^z��S�w���;N�=t�O�rZ�)����]��*��bd\:ܻV���n(4���c�Nh�Խ� �$�o�yj⚑���K�yW�y���N܃Iaz^;�lݟ*W�4W׸?<�0j:�5�߶�n?��5��٩B���T��aQv�׀��tK�H
(����H3t� 9 H�t#!ݝC(!9t���Q��w��0�u�>�����k����Xt��z\j����b�_t"6����^w��>5ol���t[_%3�1�u6�B�P���А�����x�g�y��%��^��<��{P{��T��C�v˱�V��Q}��q>���\������F*� ��� }E$�#^� I]�D;�:
qǨ�'/�&�����^s�жZ�J��.-k��
�D=���_� �{���:G��c�����/��Rw(3zg��OQ�c�kl��}Đu�������ץ:�`�#�W�!}��.�hHD_�6\Q������ƨU���i<
oK�rkk6:���N�'>�K�z(�)d¹��G������ss��[l755;�x翡���p����5 `{k��x�ި0�gz"d����S�D�5N�9Ws�A����g=�D��I ~e;H�C�y�@ȵq��Ϯ�f�Tx��ZR�Q�{�:/�;(��U8x&i��&�`�`�u�Xஸ?Y��bLjP���V���_iN3��r�>/����k��~CÜ+l�U0�y��x����n��E�y��&�[G^E�Ƙ����ۘ�0�!D��m�^����{c)������2E΋/36I�)Қ�O���3x��+0H�B>��|��oH5�Lv�'�Y�G�-��w���#:&�5�ˈ����Ɩ�C%�[u8��B~�[��xW����AF�f�H��%t�(�@�amd�p�z��Q�p��Nm����������mj��˦4¥S�B��:�n�������%����$���U՟. a_,33��:q�G����c���ꗘ(�x�_9j�F���Z��+5R�U5���� �@U���6��k�cUr#�,1v�fEd�]�RM��Mxv�BZB�]�_�o��	u(�����J��>G����n|.���_�+
F4\�exa2�)��
��M����~���ֈ}�fϞ�
����%r���~��e��?=�Wn��%yմ���=�^b�uF�-��c�pѷ���#;j�!j-��t�m���%a�D,�:�Vv���T��#��b�.y,�0����qu��{��(�?EУ��4R��:��������ߪ���@���0:Wvl��yf�~����i�")�� h�}�b��3�M���
�=(h�:XV���F�����$�Z�*6�,��`/V՟d�
�+0�p.*�N�Iu�8A�]�ԿK}�IU���Q.:��}��������{8�|���nѦ8$��X~���E�������u�/[C�<�5��m�5��]�к�����
�꩒@o���`V!��0}�!��������u�Iª�T�j�* F��,��%�dHEɛaEH���U>z	�!.ׁ��8}v�q�s�:���\��+��hi�b�$�KvR��52w#	�RQ��>9���Qy����%��=J�i���������LB5��¥xԝ�iJ[�MC�
vo�S����|:��

b���鮜�@�f����G/��j.�����5�P��=����I����e���^���i�����@��d�,��D�5��8��H/�C�c�K+d�"4�y,qʉeA�·���](�&��X2O��I`B��8Q)�܏��O����U�:'c8���	��L�||>�[����p��Nw��S�.�BuH��쑲���c�:?�=� *j�����$��\��O �d,/!F���]<e���C{�KZ�eCܸ��x
�C�g�{ e��?����Q�"��Х]Có��w.�J*���/X�{����H���}��!�o��gH�<�Ӗ@zܧ�׀��dn�^�ϝl���4��@�&"��� y�X��`)79ͥ�띶Kf�a���Z��L@���wU�Q�G|���N�u��v�L��lD�Λ�w0o�y���:u�U瑙���R|㓼B�C��Y�h���<^j��I��:-y��� s3�U])/����*˽��.����h��@}�k�sjs}�E�/w�P���7�Cx���U�Z�h֩�r�8P�_S���{Z��F�#�R��^��b6 �F���*�?��M�DV��1O/-N`?�2	(��s���7P�ϛ� ��n�Y��<��j���=�/���#���|(N�����%yD���I]��#���ભTδA
��Xuh�Q��;��
��?6v��\ܙ�G�Ǹ �E%qDݛ��6�KI!��RO�~�o66G��+-�j�BSˊ�s�6g��]^�>�֡�XH�:��U��G������'|�"ȷ�[��Y��-�����7Xf�\0k�[�m�0��c�$���=���O��L�<�K�e��9՚'����6��k� ��~
�I;C��ڥ����^��unHT����9�fJW$����C����k�Ul�Ȯ=�����獝Ǻ��Ĝ�R���������xa�m|+��>��2�l>�6�X���V�cg��_���k��e�R�X}��]}?��J>��Ǐ���}�EkJ?)�Ia:'��c���I`�2����z�R�B����}d�c�<�D�"���_q�<����~˓�"���͈ܳ���<�bQ����
�>Tuw8�w���v>(�:.:�~m��w��|�jZ��Ag���t�`�-���w�75��.@Ve[�")����X�ݱ��$��3�-�gB����)���jEy�D�G�v����W"4-�[)��b������vI��)�a|/�jj�]�#�F�/�nM߷�<�(�ț�qH��:�ѐ����0��.֨jR�UZn�g0#�q֠�O�����1�0@�o��J�+�\{��G�QS��"O`bz&6��+u� ��s���Z�L�KHR/ Gg����K4�an�����O3oq���202;�</�A�ǣl^�<�;ꖺ򃧇N,*�W��O�����`��iޢw�y	,��(���3�i���>~�G���
C�2�������H��e�Az�K�.}Cv��x¥c/�˨	8çb���]@��FI�92�.s�C~a�V$R��bf�5;��K&NSZ �ſ{�M,�\$u���*������m����fՠ#�4�|^jm������m���ׂnK��`B%�VV?D�ٳ�ҩ����=���֝|���'�u� ��o��g��N�Lx�(��*铍��f�;�Z7�U��0$�7L�^O ��f�&)�e�;x� ���5t��wI�d����ㆼ b�_h����Ej�4�˪��� <H��OGLn��_�p�闁��(�0�4���"ϲ�t��5�#lM>�zf��E̖6�$/���;�����kt��
|��C�!���������y�Ă-H����qıҚjQ�g7���cA�p	D2De1�|c�R�L�(��W�~�~�\�� v9I��(��w;�R��[OFTնk	9�.1<5��`�,r:�}�MA5߻s�>̘��B�"aߏ�)��P�Rտ��)3��?B��y�	z�{��%��`"�I���jg"�JCy�G%�dB�R�Ƚѐ^���j�Ma)�2�щ��$���Djm�ѭ�P��(ʺ�d6��%_�r,-��y���Gi3�q��=Â��kF|I@w;CO졏�b+��D>f�)L�� 8���#%s��'��oX}\�@�ET�'�?����>��ἊSKQs�K���}9�ɘЄh*���]E
՘
9ەt˸�I4�s�GZ%x�-�[�x�y�e���4H\H�o�~�#>� �&l.��˧8�}D��Qޖ���my�ǥ�J�`[��{	��J�Ӎ��0�ˎȤM��Ӂ��b(r�k!y����z6
՞�Tܺ�������/U-�1�]I�#>�=4ʭՙ U|.������@>I՘�E��°Gl������}�e���5-5���@ԥ8�e�w�m
���D�o5��G~S�qzފj��^��L#����}�bǌJ��4��$?�ټ叾Q�x��4�^�}ފ(I��oTE�~ƺ\A*��]�=���3�|e[�yM/��Z15T�N.pW�Ą���G�l���y������Y<\�X����f�T���&D(��s��ǃ�f��|�Je/=N��~#S��PDȎ��8�?<q"���%H���1������z*I�.�/eP�;�MY����#�A�q�yW�:}���M�ճҢ�����®��(�fiy�\JiE@�j��ogw���WG�G �\�K��;I|p?y� k��դ�f\aKރ�4	������_<з����?M����6���/xN���z�n��wD�f�@�h0-2_�C�w"~�&��Om&*�h�N�ECa_>��N����_,�6�svw��/��
 �︨���/}�(�-�P�#ܤ/�D�O���j��,�J[�>Y�X�-�D����*xT�@:�I����f�SU��:I��>{�vI���s;qx�W���b����-b%Y��2���^}�{Z����NC^�⋢�c~���|Ul4�+�[�x�3y�,�?�w�~��q͢i��g02YW��R�W�u�U�ݭ��w���EӶ�y���o��h�ˏ>�Gj{����pk�ƞ\0!sI�C��a��o��"B�`B�8tĥ�p���9����׹Q�����zKx���
o�WSQ���7�Ɔ�5�!g,�3F��!��2��͕�A�Ջ��F^����e�V��^P�L��n��F��
]�Zx.3bza		�w0����.��t���O�.�E��	���)ٓ�pm{r7�3Qe/2c4ur]�Y.R��[䄲��������'�ϱ_�_���/���a�=[gX�}�/�(UӺg����84B��� �r����0?�d`�P�Ӝ��
��2fq��Q��/���\w$!3t��@�<�o�[wXZ��i%<��%.e�<U�ZK�W}�ϲ�:whO���Na�H}'�2�.nx���y��g�BE��hi����/��h��@���^��(C���s��4wkG6�h�i.�h$3�ES��=���Z��-��G�iIN�N�Kzf�����s|w��������/&y��R�G���Q����wK�X��g����H9#��{�xv{K�x)�����̢��z���jH�C!�a��w<��Ҕ�Ul2�ژT�b��C����!{8]�:���CfK���R����8$lx�\䴺.���*S�c�v3ٵ#9�)m~�.�㑒�����¾��˅������y��/�������u�M�{��(j��}ͱ�BR�{h�N3�DQH,����=)�����i�gql�fa�N4��T>���q9�=刵$��Pb!���gT*�H�y9O�����w��F�|�������h�ږ����ުӊ��@��nf<��d��8�]T�G3���Ҙ*���1R�ti�����5�P{�J��{��L���gd%�bg<��Ə@z��Vov�����6�5���	�wG�c�\�/��H�ܐ�V-��k9���ʈ弓P%Z�k�*'C
���0��To�!|�)5��z��ċ�
8?��F�7�ahu�o�a��s|��������"J�p���{�iRKLQ��Q0�>Sm�yN��Bރ�%��j'=P�޶�7�f��b:�uq��E�;�|FT������wcJA�?��z���|1��	](�Jl�rx)��N�.�?��j})��b�}�l��f������'�N<%r�s�z�'Y���Z�.:� ��P���)x� ,o`��9H#Z�F`׻"���r�y� ��kr��E�D���O�g,�Dc4IYF꺜��~B�{�hθ"��m-ݻJ@U�'�!ң�_=��@f��e4�Z�R�¾�e	�}N�	����R>�0��}�N�k�eI�u�9}������_�G����u�U�o�æ3ō]�$��N����A��q$�$�
�R)�ENj<L*<�6�Id��fVM>E�#�������w6I��O�͉}�b�J�ɦv�
�	�dx'���3�׿a��u��n���6�z��;̙�ϖ�5���B�C�+]�:wW�~����L:�c�ż2�qe`>�`��������y!?���gv��(��P��oO�>[���P���y���Am�$׍�ۙi����V��h�j,f�B�ё}��K��xC �eǆ���A�����n^�:��> �F��x���n��ŕ��H���ۂ�q�oʋ��sQ��c�z�����wu��-[��g�ªT:0������[�17)o�ͦ�9=Hȑ�u��g���\H���������{}R���Eۻ�l�)��Қd�$�9�Ж�n�>i;�W�<�������	�
m�m���	���n@��Ė��9UIy���%���(Ր�g��
���n��/�f#JJ�L��i�����G}����b�4K�WWW_��o��X�٭���A�Ȣ���Բ�}C���ܿ�r���o;�� h��Ѹ�w)��~��t�m�s��y!I���I�d�=w�4-
l)��� {n�c��)����}�1��o���cki���2��+���L�$w*���M8�}���@c@��v���Oh���:�ռ�?ɄC�M�5mp����bJZ��c�q7Тc��;�wUOV�1'� ��ήm�~�@�1UA����[�Ǒg
nZ��3%�|SxD�>E�Y%�{^��+
9�fR��0!�ª���}xxx~�ױ^��~nj�oIff��Ű.62�'�ǿ�����������^�����˵�|�-W�"�}�9�F�6NZ	�~�۬;p��MF���BAy�Pc}N^ڊ=�^s�u,)��iXL��1�?e�
�m.Jr�������d�9֞R�L�]�قFBK.�iF\tb��9�<�u���,�Qñ3�ɦ�i�cI��"-Ɵ���~���]x�@BA��F����U8Sȋ�WR��7P=M��{��;���[E/ɢ��x/�\��Sҗ5|�����T|�ܽל�fTZ⻓1�;�O�V�:��P	ucb')@hW�ש�����CzMD9I��w�[���#KEBT�»�C@��>NnFa�%�Jx�A���E��ѷ�zzQ���|�ͥ�)�8�5$�`A�`�D-�\2��)!?����m��K�]e>$EGo�r��$���Ml��"��J-��Ը7pDVʴM�ӛG��!����J�0�s��AN5���bCR�����Ql"~��KfRm&#s�.�\�ȃؾNb��ι��-�����ٓ�q�w��4��~e찺��"�=#�b�f�a\���3-��\��}6������/(+�TE�b��Dn�.������c�:[xLZZ���Ni�g6��/_����M�.������h%�����]q�����R��~�j��o��灔���$�8�!�i�9�i�]V_��~��"|�� ��:D�aeqYz��,�G��jZ:����]��q���K��>��Qag�� v��tㄟم.M�3�|$S0ImR;�xl��o�б�ow|��z<�7iU�����a��Z��g/�˵B����NM�ѓ���&E
W�<�ŉ����޳,ˊ����[��|g�A����k�����5.�dwc�Wg%껲�F�W��� �d���Wsa~0��� ��Y�lW�H�����o��*k.��(-\C�0���5��Ԯbo����K�޽�!n������+!��Q���5����2��-��W�@Z��i$����,�X�R&Gb�w��tQ�����r���l����b$~�e�c��VΝ}9%�����L6*Y޲RD6�� �r\�Ԍ�klޝ�����3��92�7[���6��H�4��o�#($���~�����F�vYYYQ�U�������_=�v�'"�-�}]� }vi�Ŕ�>ʹ�ǡ�'������)7b�fb���7�r�tఎ�M�p�^�D�i�}�:J2�r��'Z�{6�7I�&Uo�8��B(?7�X�0's�cN3'�U5"t̫h��~��AS�	ݷ����8��F�J�[�"�[裤���~������~��v�W�G�c9��A&��+�L����v���n(���u�[��*�x�Nf�$�?��E�ҺAKk�(�0)ro�V3gk�����F��zo8�=I6�L�wM*E��f}��^���j��[�]&w!@��nC��r~��|��[(���*�Bn�[���Җߧ��+=,�F�ܞצlI��XǰChZD˃	����23p#G��\���e�xp"�m�jx�j��M����K*�υ<Ag^ї��4�"��i�@���e�;��Y���:��w4��r����%D+���=.i���Ì���u�̎C��X���:���@n�Rh$�1����;�Z��w�gB�K��փ��%�:b!�%	˼�>9����A� x�>x?��Y�]{�����O�R��ly�
RH��c�!Z�$���SC��*\�_���q/�lD%#�O�k%�O!R�\ ��sF�2�֛>@ɠ_������='�0�/V�E��%�֑�������_��=��FQi����o��YP� ��?����12toc�zq��k��iV��薬ے��fz�I�y�t��O�=�����NG<��[e]���Y�W�|[�E�N/<�n�)qW'8�_��1����;sBP;b].O��u�JR[��*;���m��صDX(|�h�8�rjl�}
<�!��_d�w�ŷ9��_�ߨ����W�>�گ\�� d���T��k�O5zNj�-a�΃�N�Tŷ@$t�-��H;����l�zC^��C���!ma��lnԚYl�!�|)��R���Ξ~k�}`yR���+A�d�G�֟����	;�	��M���JBԜUw�#v�Z�2B�/�z�[vG�e�[�K*��;��q����O5k�-�{�fid����ʴ��hДgF�,$�S���mS��h��E�8ʤ��i����f�?�?�,]�V�߲`D~,�����p��w���n�74�I�����?�[���g)�tZ"�M<g>-͗���*s,X�s $�k�������m���_P-��o�m�GW���i��@���A��qA���!��.��~B�
��y�N�e������I"$�S�="�
u�!�O{���M�ȩj{��4��f��sJ5�wg�HG~m$�յ$̬�T��&��c���Z/8���lq��e%9:�h���[�M�d����O������|Ugx�<`u�)�O�>��y~���m?��4�����l�R���JĴ�~����]�J"��X�l�J�nx�m��/ 8�7<(|���u�;m�q�nQ�)��vX�ܫF.|<�)F�<K߾���g���
b]�-JV7���x������D��W^v?��<5&2�Oc���E���;!����u�>���i���p�D��V��Lϙ�Z?&��|h/�Ճ�Vf'ڰ��S~%&θ�
ёIΓ��Ť���+N��]�B�r��|%��Zi���J�@�j�ҩ�qkn��ZL%Y����N��`���i3���)�J�^��@����f�Ebv4��fL�@e���8ٛ�u"���Y�[Y�ݦг�R�/�_�C�Q�'�ݖ�����@t��Ϝ���n�j�g,X� �_	���6�j%GҾ�Ļ��J�v�s��~d�de�6<�Cr��=f��c#i������wY��tf��~�.��ɀ��UNd��m�H�`�y�|�7����t�o�Do<�H�����^OW���'��^j|ɶ��W4���ATu$�2�.��;U��y��,Ya�-���1?�ˋ[	�����&��Fz�o�0Ku���y����m��J������;�(Y��T��~�v�q�%;o��w��Nt��G��?�HD�>�wK�i��@�^dw�.URQ�y�eb������HY�n!>q{cՍ��\T{9�]jS�R�G�9U[P��\Zz��]?F,ۏ�GX�]���٣��g��Oخ�̎|�:��Z2��b�e�on=�\�S�/�N,��u̕��巻�]���a��gI8�"�6ꄮ�j������<�\��Gk\��B���fq�U㆚>�٥/.�_����iХP�pT�&��-�,8Y�c�!E�����Rf��= �;����qp��TO�
Sݦ#!9��і(�M���^nDtBfz(��Y�e;�2bW�N>�s�����y�0��ة�w�:@�y�:����9ʮ!�p�]rM`4�	�-Tۆ׽����(6�U5c�_S����B��/si���>��r��o���(��$M��8M�h�v���mVoa-����(>��XA7�	�6D8i��W �W{�e����v8�|ǿ��<�R���كL$n�i��nh<.�:N�R��Tb{�eM&:�c~�c�Y���׷�4aS�ꅄ��¥_E���Fş���#ABz�1���&E���3Ya� �i�A���\N�MgF�m��R]l���[�R3l?R.�1���r; �b}��oI�yFC���?����{3 ��\[Y���Nw7e�W�� 
[�۠�<��xi�w������j��ۦRB���	�q�̬n�
�����%r�p�ћ�Y��5�|Hd?���
�vjn'�	�i,i�^��ỉ��Z89�4z>�[�>Y�H��p#!�Gc��158>-ĵ+�0��-CFB��rNzL��|�k9)aJTL��(|����a�h4ۡL��x�r&�|%�溹T�">����Ƨ�RSQ��TTZ��~�8@�,h��F�l�jT.�		�ӹ�K�_�l�@�a��{����WCB�$�~J�V3�KX� tb�g���rNԡㅸ݊�9^��bx
v�]�=�ee3�@��٬uR�j��\�f̫��� xugy�<�!���_��� �h}#Ѧ/P0'�<xt�)x�I��V�-^F_������4��aCB���P9;��,��0?_n/ٽFmߐL.�?��5�r��;����r�7��f�B�Z\������䪢JIr��jlO0'm=��*8Yq�VW�/�>���J�q�t�w0<(�YodV��̻:�}�*ў$��[�:�YX��ܐ��/��t/*��&��Lx9����zM�|4�dN���h���B��ĥ�oa�#�Y����k�Ǖ���'��|N.O.���]�KR;y��|{5l�z?�x�Z�����n������$U��&�iq!���3v-#[	t��tu���C�D&2�Ճ�<g�.#�y1�i���I��L8�I�־&m�����ݜC�DN���*�z�X���s���\�8r��x�B��� �`���|��ȵ����r�������:��z��!��Z;P�c�;�q�~(Mg�c��ZFᷟc�kh���J�<�'HH9Y���Q8&�-WkPcXee8�W`�=Ԏbj�n㷙�T'�j)IXH0w�
Y����i��� d~�$�j��6�:�KW �y�#i�Ey�&��#�방��&Zm-��\M��������^%�o�9�����[�57������$��^�La�)��J��;��EJ����ȊH�K��~H�f���b�(�۶�*�����v���ULdF"����1�Q0m#�2T�"�\���@ʢ����x=�t��v�FF��Á;���[��a����f���K)�C��1�?��	Ve�n�Y������|�q6A8�d��S?�)��d�5�xXŧ�:�S��ȫ�#�4�5�d��)_����)K��xC.�$�r�3��S���q�*E�j:�/ZJ5�.1uA���W�;2�`�) ~��Z�p8��'�U%�����Kf[],�w�n�s�]ƛ%�a+ku>};e������@���)�|'&E�� V��h��w�;x5��k-|�V�݅w�"�
�M�R��b���w�:��Y:�/��?Ўe��&CS�����2f�����Ζ��i>�Tk�?�_�����M.�}8��y��c#6_�P��}8�]�=� fѐ�%����ګ�zgw.6�
�� ׍-xc�jղ�T��W�n�(�LY��;C��ܽ��G��"�R`�b�^�ՂKk'�ԭ�[�]e�:�&��S���v���������׮�L�Ԟ���QK��N����+��*;�T7���MB���mm�2Pi��"$�K���Y4�hm(Ť6��nlY#|�Eft�����a����Z���H2	��Ԭ<��V�E���Cʷ�
��[���oeׯC
��*U�b�X�(�f���w
%<ǀ�#%0��'��gZ�����'�)�`^�<TSW�b��yr��&m�&�.����՛����S_���R���"��y�ȼ��⺾�G�9M���b�i�����O�翩Q}N2M̆�� �: ���&��uem�A�r�.��A�!�1��"��`�T]g��#�܁�	���Ce� ���i��$�� ��x�yg�W��ũ޲��e_aI[y���b���K���[�xgl+��n�qV�т�kx�ʺ��I�:s�еC�!��x
�4�K��x_�n�]�6�VU��k�a2o�:_�v� ̽ˤԛ1ki�WϢ�K4 ��Eؽw�E�>c�J��4)��p���c���s���k5e���E8$!��J�m�bX�kIZ�_�0={VWg��d���^�ݨ��%'��K7N�MG�&c�:�@_����<��E�'G������-�[��}�ɩZ����A����/�0�T�Py�f9��E���c��Kp͂{��+����{��z�� �p�[�uf���]�ЌQX��-k�K�OK�
�������I�q��mf����=tsZ�ҝR����m����Z1
 0���ȨPQU$$4��� ��A�&F���H��!���n��C���9<��3[W�+��-+`飯��X6CT�F���h�>|v�=)���x�;�C�������(��Z���4��c�3n������|l�!�;��lu�&��b[�e�5��;��$��tq��Yɫ�o���Д�o�5wc��	|�:�A��� �F�n�,�P�����w5w�T5�濺K��T���<��S�O���Jꠘ~>�:�էo���}5���ֽ��k;h�t�����G�r��uʴ������ez�������f��4��	���u4���1��)#��\�^:���t-���ܬAO	L38@���m�*����{y}�����ǆ�Ӑ�!�*�E�M)��A�(�����k��� �s�C�w����&�|S�$H��M�x韑�f�4��gi����p5v��,.~aޘ>�av���Csel���[�u�2��<� Q��<��b����ȕ��%g�=\IFW��w8`) h�ӍD��#���YP7�^�2�z�SY�Y5���5͖~t��TH�p���oI��>�K��m�������ԧF�(GT�Y��;����.;Ti�y�֗�N5�k~�גuQs�m�݊�=��m�Ե�|���<���gх7k�|s�eq8D���'�k�B:eT��z�1��KT�<��Q�����?S���ki�
k��ReE�@˰�շ[�W-��B����Z}�ε�p�G��1r��l@�$[����M�k�.&w%!9I���kP �ӿSjθ�g�����M��_�Ez8%��L�� �x�����LM: �{��E!UI�2�&B@Rl�%�"p(=y���ܻ|A��kI�i�g߸h�F��ǺN36m�����F�p����(��qX&��#+���\Uq�a�Qw�f��Cm�1/��#p*���{q�(��p�����dC�c��V�xW��6h%��!�+x��~9}�s�e7�2��d4R�vPF�tq��]|Lr���g;�=�6�ރ�Vy�-�G}���WDVTҗ�x~�[��f�l4_��q�[�]���/^�?]3��D�K�,�xM��椆��y���t^�����{�Q�we_�1�@�ql���2Z��>�<r��L��Z�����N��8��r7�4�Hp8�qy�^���7��1��^�����V�����G$����Ԯ�bE�Fl���.����)�I����T-fnM�xx���_ 舭�JL�]���.H�:`�	�A�IH {�!���}-[]+}��	c�S�����v%B�� f�5c
��ܛ�(d���l��%��4��;������an}-�3�mp3�0�J���x������!v`�3 ��/?��e�������?��9�!�޿gh���}���||��h�<���?%��D�PK   ۍ�X����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK   ۍ�X�ĩ�xa  na  /   images/c9c0af01-d4ea-463a-b9af-0ddeafc58269.png C@���PNG

   IHDR   d   �   �oƬ   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  `�IDATx��}|�����ӝz�\d�Wl�ml��!����蝄�nB=		=�б��ٸ��-ےe���m���=�I�fɆ�?�gI{[޾yӾoތ�PSU?���ǆC��_�;��OHQ�^��#����k�G�X;�����V��hQ�c;�=X��� ��c�v��?�����;1^��d������(?eohd��A.��%�9�?;� Mރ�!xI;̫V��VZZ:pԨQѼ�<Scc�����+-�����LxF��9���jZZ~W�������s�T�`��T�_�����S<���P]]��~�-��۝b�X�Vr8�����}��%���5K�a�����N�M[����4�����t���oG��f�q��l6[J��������w/�X��frgܞn����٤�-��C$�m�y�~�8�q�ܠ�}�O�(m���8����:��
�e� ���s��Ü5�|�j�?|����ZŅ�s�y���͵L(�h4*���܃�ᣋ���ñP������{�#��7�s�u�!������_Uͳ��!���4l��XC]�SO:i��{��nQ#�ǭ�Ǒ����w��HE��]I��똔�I;��ъrRxPc�dr�S�l���G��2���(
�\��Dh۶mT^^N�~�)͜9�\.���4�����Ӛ5kh�ԩ]1hР����.AZ�������Cٵ�@�����G�����}�q����7�@*�WQ�vf��m� �	S(�?Qx�f�HǗ�C\�\H��A���y��`��4׭�8������gC>&> ��͛i����EpDCC͞=�����p~BL"L8&���ٺ���R�����Ea4"�0�/!Sv�^/O��kn&�n�*aDDZǟJ�ߒ����3Y���z>���a6���59�9���v�����t�;(�
b<
��ʔ���DL���?�G�'�|����d0��p�^x��̙C�{�<�Ν;iذa	g*�_�/�h�/?��ןj�aj�m1,Ń(�;�>�(�*�[�l'��~������jӅf��Ԡ��<c������~d�%�8� ��ҍ�][��Hq�;W7�M�YZ�~�_�	��N��¯����۷S����EE':8N<�\�RG�29�yQ|������%9�=���<��a�q˽d�<�n�Vƭ#��ߙdP�?�Y�g �0�̱d�5Yh`}�T�6�H�\:dM��R�DW�j���dee��2�А!C���9;c�Z�n]�q�$|�$�Rv�}b�"�|y�����I�>mH���O������~�5�L^��x��V���T%u�kv�<& �`��Q|233i����k�.���tҭ��J�����݆g������$\a�H4��k�A$٧K��"
�ZB�_\��Fs�yy^{�bU�:]B���^wsH4I��a��I~�t*D��S)���H�y�M<BײE�B��ޏj���l�FX�F��s�)*��n�����pG�� �F�I˖-��!��I4�(P��/��ig�x�� �_^J�	��u�!-�ᾭD�)#�,��)�w�f t�Zl9���l�)�f:��)�<C��-�Mb�ׯ��w_Q桹�y��0���q�����iI�`�@�HO�ie=�v�yV7d�ƉLg}5���%�i��Xd���:f|�pӓ��8d��(Y��暮8�2z�>�>�5���d�Ÿ�ފ�W����%a�[���� ry<5�{3Ew�9ݚ(<ȡ47�<�TR1C�YުJ����X�-o|��/�Y1iy�4W���k�PFَ����XL���&�NQEM��G��$5 �����V�E�y_u�G�"KD���R�1t8.��x���]�+����G�#snEvnc.I��|�I�*����9H�Y��Z!�:҇�����q�U{)��.8�v�6Wd\sEJ�Qp���i����.?���EU�=;)���O��Vi^5��|��K��I�5���֍;��&��g
QҺJO�a4�쒒0��S����Do�Ĳ^�;�1�R�_���tw:�<�Oj��&�}�;���V�%�x�_u�X���cRYx��?%�Y�y�	M&�\V���K!��ځ��Y����kbH���VVo��P�&�.�I�R7E�蝮G;6 �K����X����CR���*������3￞M��X��|.�}��;o�n��|�Y�M��������+�7L��)8fL�y�� �����'8�>a�>|�Xp t"��an����b^�(u3;r�.z��X�D�vQ�?!�1�x�K3O�*"�b�f�|����+`�ܰ+NR�X:�k�&&�\0Jq�"D������X��P���mC�Lj�׹ߔd�w��[�)���:D-8�ȒN�Z�>�	O��1�~t.U_t�EU4q �$�y���	g��_{�b8�h��a������5E����3�>Ņ!��*�Rc^�(�̺*,�$�?�,܃�b������4q�ZD����2e�-~��j@aV(��>��V���TX^I�MM!�O3���-�����������鐅��Oپ67�1@�[,����r��B�R��{5��G!�6;D����(�1
{���\�����z�!�ȱd�q,�C�[��4�=|�4Z��	2�Մ�+[ D#Vm�!k�%G�@D5�eӒ�0������6ԏ���d�i�Shڧ�)����Sx0asB	-������Q������W:���r! "��ҵX��x�TQټw��r�|��YbP|=����/��'\5�x�K7Ӳc���<���}��n>��I=�9%m��q�A*]�5i�뎡B�cO�i���L�����~Vu�t�)L�W�vk�&>���k�|��h�Sx�Rr��(5�z�̐6D�\ugl/Њ����Qp��4H� ����X��X��g��Si+�p�p�'���'�{o�ZQN�G����^�������wʿ>�y��|��#�hW9���N��J~f���\C�<�{w��%�z�qC��ɺ��d����a�;J�����M���C9O�L���QRR�29��b|�����1(_,"aU(-�[{�@���zA{��o�7�ob�i~�j@��=�,^z����w�{�H����E��x~΢�H�3��i΍���L����R˺�x�8�X����ȡp�ƾ��� ��iT����j�(+,pt�,s�n#SV6��6�1�ؾ
�ٕ�ʌU������<p[�n�ݻvѼﾣ�{,�c�&�1�N���+V��U��c��t6�G�)���ϗ~+�!7�j��}��)'��d[�����yL1�<�8���-�q��<���|���v&=҂>X�V�1�	&�p�y���E�l�k4u�\0T&��5��^b����q;_;Ơ�`��?��h�B�5�Ӗ����Qf�3�ƃ�}G)���+d�����^�E'��F�j�]�'ӡ��SQa����b���\�����%�HXL��5��� Y$ˠa�oEW,!�i3D�XǸZ�a�.�'s?sI�.�B�'6l�f/e�5�G1������ٿ�n�o�@�f��E�U�@�&ŀ��@?�οX`����)��N~ha뜇��2zxv���_{�u�}�@�Cy�z�(���)�u��]�5��\g6�l:�[K^�yi�TlRiBS5}��5�;_��G6�W�h�%Bc�3�/� gj̠���/���%%d��>�!�Yoe%�Q͔�*ں1g�j�%.+���ɚ�My{*e<y�͓�ݦ��w�OX�;��3f�ʍɝ�FR���YY���l�Ŭ#�@�� ͑ȧ������X:7���M!�`�8�M��&�����q�]�����(p�*���V�������x`��I�WF�e�*;0�?�][�6�E�n��Q�:- W�iM��Jg��6U�U+.ؘ���a��rr)�JQ_RW��~a����TW�zaIX�VTF����?!ӐaT�f)�+���x�}���`�Lc��?h�f��$�N�}v�q�k�?|,�l�l�;_��/ba13j�귣<�A�E�b�aג�S���6F��/�p߭dz�~�-�c�G��Qf�ڎEMq��e�Tߵ�~�j����3e]Fc�E�	������>���Yw� O��=B��K��D���RZq�Dj�J7�b�)�7t'&���;i������eІ�SUG��ScN�t�l��ݔ]U��Sq�{��NVR�[������l�2�Kr2����v�`sT��hb����t!|l�"aa�9�=�B��Qx�Z��WC3f͕��=�4�����>�����!�$��ffm��n|�3P�51���7���n��4�9)Y[��My^T�O�q�S�u�f`W��97_|��*U"�o��zX����G������=�?@#VnbU�-�t�=$��� %���&jig��]*�x�a��Y`�����#�t�ƌ�G"�b�
�,�YΆ%Y�`݂�)�E7y��l�/��i��	Q�Y�����Yh�r2İ8��d�0�� ��A{��Iʎ���=���H���k5֗�?� �"���BnM|�5�A}X���kɲr1h�AX�?+��y�e�XY^.���a&s *�ϱ���4b��Ɗ;��P�۵g�{��%��JiJ�����6ho�n��Ԑ�%�2Y���{�3�@���k��Rz����i����J]N�mٺ����<�rʛ:�|��+I(x�⬫�pG���W��cH��&������"�f= ����#S������N���B�U�x��Rr�W��
���J*����5}�	��4��	���7Ɗ'��L;�r���ތ�F�`5�WTu�r�H1��r\.*�̤��f�()|Uߛ���N,����gb��k�'�R$D�ywf�$@ ,�bXeeeǏ�g�-*";_��x[(���ส�2psiZ=m<�+.J����W�k��G{s3i��S)�tp	{}<f�2�9[�nڧ�Q6~'8����::}!���J�=ӏ�̙O��Ĵ�ef�����jz�vW7����8��*θu������xa<�9ܔ�GYz�	R@����x���{i�1���_��n��Y�wX�a�c�bDI��m�0J(jG��X���淕hLm���1_�2�$c�a�i��ZzɝQC�f5�l�<P\�T��)��`{ �L-;)OE,Ժ����� ����/���� ^J"`,]��j E�e�ыx��+ϧ�G�%Ǩq��aw�<����^��i���E��/���6:R�_pL�P1�;�3����4 �||�+�!o��\�^�-#F�)3�����g(��
2��e���{s'/�ba��@0(�:5���}&hMf�>�P/k�x �w(�0+�3�&S����= j�E�
�8�ڻ�7A�+-� 8��c������(+��%}��Kvo5�Di;�,]V�#�˘ �n���O>ok�����o��虱X�-�^�N�4w�����p�P�B|���^-�(�מ�؇oR&�S�zMQ"���`�.����g/�lV��������c��c`�`J#��5��BU4����v�k�>���[�Ą��z��am���X)D0�qa�cT��Hٶ�����}= ��!��w��k+S0-�@{���{X�!q �[�x2�@{��S���d�w0_<�lh1{�^jWI%�G���-�O�ٿ�t���AZD6��O�'w`ᬏ���\��~�__ R������Q��O?>�-C��컷K8�kL,ˮm�nYON�#�i�-,���	�S,���/ܵ�B�֒܄�C=z$�a-���E��/"�K���d8�@{�@��=A�d���%	��|�N�7k09fڂA�;���DX�RL��@s��V��a��.�4���ŕG���C�~2���"s�df;=��KQ6}�6+����;��a��,������kv;DƱ���i?>�p(�~A��[�m����$�|Lm�.��v���s�4z���A��>+�
�a0{��s�I3�1q�;�g4l���3����`�5�a���KD:N�1��Ρ��}T����XCᷚ�3fA���T�� �!�PD�ē�^���T�f���3�c�9�#t��q+��C�la	k�N��4Q�Z<�dYA��FR�ˊ�Ov\@���Հa��A+e�ב��{��j^��7,/�P;��WYX��i'�N���O�dE��]�E�{��fn��b�N:�TJ�8��K���k����~,���J�2d�,TEY\�[C{F���3�]�Y�����ߑ<���{/�T*~^�ժ��f�Y��6L}����bmo�"zd��4`{Y���"30C�]M��J�e,�G���cy�+MvSur�(��i�y�q$}�D�&���md~�k��=�soH�7���u������dXyJ�y�\;+�lW����f�z���ࢹd�q<���"�g��o�Ҋ#'��2���O�`;z����E�$���T�����QB�v
�h��]����������(�a�ch��23anR�ih x"���5c�ƗLU��}~��
z�^����2�����*	���|+W����i(������y�Fg�� a��~u�@�Pd�z6��WӌY��x".+��w�z�Ǔ�hg�(�N�^;~u�SU�8��@�F{u�����5�D�UW��_D��6����-40�&a����4i�4���,��`-{˨~�zY�u�������{�z��/���hn��E�6�$���(�_(54��5�Ll� �%:��o����g
 ������x�ۨ��W���׮��7���㗵$��������E��BI����䌶7{���@A��w�t�����+dcΕS�Rp��2�i����<�g2��e(��;A}}ͥd[��,�\.���Ymϡg�>������|/!F�6:���rrm�v���e3�I##�h8<olCÎ0Y&��O�K�+�� >�\Ua�HEE�wj{c��"*�@�����h�D�t�8�d��T;�R�d#�I��y�H�LBVW?�|�W�M�A��Ǔ�SI���ke_�>K�1Ĳ��D|�%mm���(�YĎ6W�X����gis������陔�ȃd?���I�W���#���dz�L�T�փ�1��A�%���n���A��G_1$Y1̫��h���M�r���+D�8bV*p԰#%D�P3�)�Ԛk�״���O_1U��͖����2E4v~}IV\;�	�a�Xr��v@���M��ߏ.Χ���W�+�%�a��f���p5:E{����ώ8FV��%�$�&(V�)VS�f�
���$�;�_&"@P�p$�nI�Q̾�m�ϖ0�q��h����z��bS�XGK��A���Nk��%q�
ze䊍T���}��9;���N.A,*�ށ����T���b��M���W�5�		�bk���:�`����.$s�6
���^�_z�ƺ'����=^��U����u����܆�?�u��+>��(�a@��q`���lo��2.g�ѓ������bsL=��`�òj�Q��Eڠ�h�) �9	�cѫ���0V�.'���|����i���#�w�T��W�'�>�E�IV��-�q��M�8Y�Dwk� ��f�u�Z�Ym�
)�D�2�t?5@ϚI@#�� k����B� �#�;�"Q(J �e;�\�\@�/�E�[����ˡ��}��Ik0|����ؔ�9���L�Q��ֶz�B{��"�[Lj��|��X9D��7���CX��d��O�`���G�FGQ���x��Umrd�{ұ����Rđ$�w�>H���P��h����3��+(z,��0�A�ʤDFv��$���BΣO%�F�솞��~���i�9&�ڣ5j8���<OLeOE9U�Y1���Ϲ!�Ž7�=��%�%L��x�M@��$�E{mV흓�����/!���S$�:�r��1�KܾԚN��d������7���N'����H-u%M�e�p��)��l��&
-�N[��(�8����u�R�o�t�O�ɒkΦ��d��d<��:���7����� ���C���D|���A�]��t�񡁲���[i�I�1'K0.��$��p�9���S�n5�?~Or}x^�;�7�#�ȱ�8��}N[�"H�P��GG֪-� ���Ct9��:���q[ҍ�����]�eZ�h�	��ΣN&˼edV;_�h�'�-?��G-�Z��j�WL��A,�pY)�}l=f�C�@?:��!0�N;��l�Vb����6�f�u������ob�`���a��N&0�Ť�9�0r��r���)0�c�b���3Z4D�)�-�����
�Z[$J��XD���j��m�dR�.�z���L#�8o�}���j��z�d�3���fGr@p.���F|�	}���O\=�%N�۠����k���c�5*l�.2G�����g�b�еۄ��w�r�TK*��Q�\��줴K]nj��Q��x@>d)J�)!9�m�T���Ў�S� ���c�5�O�2e:!��;h��!,��،�������/<y��<�'�.ްK\�6h/q�P����+���Z�o��Q+6Ѐ�-�GPN�aX�.[H�#�&�БD�f:��g�۫3�%�6>P��rɷc����h�����j:?V'<���5�������h�a49�;ΗI�h�.�K�v��2����,����l�SO�o�>@.=u��
�)0"�Y�Y�=p��j�Kj����1��8g!"$������a?gV��^z�i����6Q�¦�7޲�Qۋ�h��o��kX�迣L��N��ܽ5���Z���`e�%_i��
�c�Ъ�Zz�v�Jt�)];����؆7��O�;/�q��C6��������R��%T۵�nB֚*M�c��c�O�X[����kh�>�FA��$���A��h�=�o�ƺ�{ �옙�. A�0����n��1���n���r
�f#IBګD�Nc�R����	�l� �����m�B�ř`y]�R���b[���cؼ�-���ךa�;'� w�&��4"��qS��F��ގ�sj��"ڐTշ���'a�X-���.�kx�X�a�3��Y�&���BUm��9(�X��r����m������ћ��C ����f/��r�i�)ڋtk�/���m�bq��5��6sQtt�%�P���KlT�7�Ȓ��E�@��R��v�j'�Ժa�� ���Kp�"�2n���MG{�bh��<^�lK��L�8��a�r�	G�/=MS<QuihoQh�	Si�'�c�hofe���$o�@���As���(8��cN%�
�}�z�(�W:��ig���H��{�M��GO�����c	����s�ϕ��8j�̅�[v���N)~_bn���^��8���W����8q>g�������tu���g�ď�9��D�I�����*q�8��~�kj����~�-���M�{$�]G{�n	E�s�<Ɠ��"a���*`[�b{]N	F@_��h��)%��/�"5����(�|.1�$^�������%�z!F�Z,�� �� �h��
d�՞A�2�lH�����U�<ST��o�n�"hoBx�����������ޖ���YL�	r�^K;o��1+���(̢�1 M��/�9������_I�a��N-��_�+�x��'؂�e��n>6��R)���^m�U?\��SC�dw�w�*���~}�dnF_������{�پ�A��:�$A|k/�e?�9&L!��2`����m��h		9�OE=.i����"����Z����8P��ʖt�� �����;�\^)��>�H
|�	��u��r�&01��r)e>ڃ�Y��l�l62��9U~��߇%��\���|�Գ���`-�.&RV;h�"V��u[%��!a�ms�;�}��q�����
���d:��V	�єK��/�u�dN�p�Q���n�"�5�U���1ɓ�*�<�$W,���9����6�#�m�D�b�(c]r,��t��M;)��>5���r�6��źb ˾��&Eljd@�bJB{�,Y�C������~�e��'Z�D⬺Ԁ�>�,u�ھ�mf�ѐgw�D����n @�fd���P���"[Ñ��y�YbmNJ߲����Vy�͸X7_$�q��E�����k:F{�"h�j����a᪘m���}�#޸3�=\��"n� 7H���ȓ}!�BfR6�*lg����/�Id�JH�I�1'��
�,P9�y�iD�F]n�{e����nX�=C_��\�Rک^��s ��͘��Q�%6 #<t��X�0�2$�6h/���cx���I��!�y5�q��f
=�(E�w�R\�Jw[�� �z����OpJ\dg�ŔG�cK'�!���m"��	2����N��5<��M��V	zn���9ʜz�z�h�)K�;e㇄��Cu	&;�%��y�h-)}GR��g�"�bKs���Z
p�W��bd�
�\�m�s$x�A\�H�Mf��-�&f��o�D��P<(��}�����ͬ�J7����Z�B�7�+�qW;djC���{���dx�@{Ѱ?�"�����7��t���^hڋ�W�醑���'z�q����׻v�x!H���>�C���r1��(?�&El� �?V>d� !�q���|=��^��;y3]���#9z�x���`I$�:�xM��;QR�q��&��Y����	�ꕧbK�a�(����&QŠ~�xF=��&���b����'�zӀ�ۢ���7M%�=[U�[�]��L�����}n�}���4���w��Vw��ʾ��4{����"���㾆`�V�����Y�X+�E9J�!���d(Ek�)����s�@�z��ޗ�(H�[��9U1��2m�<Z�& ��U5����f��bO����h���G���Nƅ� ��U��|�Xd��*��L;�~��s�,�ql�����{��f3ӟw���J��:33ɶe��������^��*1r�j�<#"����w/?����M#��&�ޯ��n������U0��f�m����Y�l8	0�\��d;�4r�{�y6 �D����	�������M �I�� ,G�Ly�O45��%fQ4�g��L��"�!���`�swh�|q�L9�D�;���řϿ#�E�j[ �����b��6h�)�U�>�0{B�u����E^�(�d[q�U7ʾoz�A펂ۨۮaw�eS{ː��{W����B�&��S4hK��a�%Va�m���\\��ؾ
j��w��`>J���l�6���Ep �˪�XB�m0a%_���b�5��3�`��0Ajq���`��ĂB���)�7^&��1�y�r���.`�ez�`N:�d-L����u����vru5P�u�3@#�t���+�>�̦�[�j���s�'���\v����7�kWSΨ�T߯p�y�P��{-06Fe�5��DʆB�B�� ���i�ѓ�%�N;�^D�Ř��#�ݰ]P�	\����h�	V-��~�l@��'�*��f!������r�;567Ӣ��!���������}��O_-K77���L�2��3>��u�5d�/�?y�"�{i�)J��B�����)}�Ggwz}�	<��JF����ޭ���E�~��2A�g꩸�z#q�UWsQI���y�������)V_���Kz��RQF{~w!ݷ������U%E��H#�d���5IN��\�l���o����v9"���j�9AJ��K�{^Jrd|�5M���V�8K�<�W+z�^�)vN��km�������7GG{a�lwc�DF ��~yŬ���������kZq�n�Kh�^؇<f+�ܺ����`�}����9it��Pu���8���/����ҭ�b[�[�cu"���W����bv�+-g���-h���;+$�2DV�h/0�P�����NXǂ�����Z?����@o������&F��A�VyiI0F�ӵr�^nR$�A��P�u�~S�Qb��t�]�+҂`�qCH��>�4��e�)a� ��A�`�.��`�PX�ơES��;�[���b�I����nWy�c�@����ab,Dȑ0s��y�>@�,;]���= ��?�Fi[>���F�n��0����Sg�m�VHl�_4�"X��@v�Jkj$�OkΣ}�QDuL��+}�:�L�Dy��i�+��j���(���.�vg��A�ZW� +��J���"��J�?9��Lw���/R��O�,O�ixzu�F�&�]L�uL{�����7�e�\�=E��)��!?;ۋ��VS��z�t���ȏϤO?{��w�eU[�0���W2��_t9���;��Ҷ�7�N&F��NwVzic0�!1�f�m&J$�N���'S��%��a�a�h*VgP;��?
)�ڠ��w�s��8�f�����!���JҊ�!����V����3~u��]D�H���?[�K-�:1��b]"�����Ĝ�a��(f&JϪ���]�t���b���� �]��H4�D��k�N���(gK,	�5�g���Wм�hİ�c�Aإ�'!������pC}�u��бl�z?|KK�a�uG3��rN1�ublbt�V����|��H��n<DaB��O����O�'�GSl�Z�n�ў����y1�ߖH�V�,��1a��D�~�X������F��\���J� �L,��AcM�/�i����e�אo��kK�3[�50Y���˶`I��ӧ��6��}^��?b$6��f��L���䑹��w�܋����"!��O'K�bj~�~*�Ui{�Uu�����z��\��f�؆� ���-�K*�c��'_8@��W�L���=�uu��0f1�
�����O?I�l:���{�L�ܱB
~�{�7�rݍ�����;�g�fb�zIU�(��(n;��D��Q�.��M���Ɯ2�̇S$��1&����;.S�{���bW���;_����aګ� �M-uRL�"�A��ݪ9��������IX�O�#ţŮ)$�t��S	����jw�bl3�>*�EbD��a��ѭL;�G��f��a�=7�9����ߑz�&ݦh�-�x���R���{�f��2��"�<-,��V,��݇j*wa��fv�?���,��K�nEA���ʰ8��،Ee�g�祿pGN�tF�����٤q�ވ���0��7��a�?f瑣�D�9M�E�ϖHNT���XJ9#�Rc�"�\k(�#'-��iNrz}7��A{[���wn'u�b7���gXƙ'312g Sp��q�8�3?d�ɤ�Y����;$(�����7AH>p i]W	�ؠ���R�$��@�yL��T��DI�_� ��ʦ�k� ���70�Ⱦrd����V+"�?c��Of����D�#��'�������*��ׇhؿ>���g���(�����$�	�}Z�`���ڻϒ*A�%a���n�QЇ��Ĩ���i��,��i&s�<�����"�jU�s��zAr��'_���.���߲�ZE�~4{s� 7y{A���j:d�jM$��E�yl�(7���3TT<��/��j*$0+��Fv�����[��к������ub�����Ĩ;��0����r/s�]Y���P��$j@{�����K�{�u	��4�6���B*��c�Hb6���'h/�2$�e����o�ꗧR���P�駰���N��(̺�������şx���1�31��Q��@��(����9�n&J��E��u�w�bm)Y���v���,��x� t~ON�&��y�쮕�q@&A��z�>{��3�01f21��GbDY�D��9��\�i�ݿt���&'L0{p �۫�U��ꛤ����h	�Xȳ�>6m=lR[~ ��p>�"t'�����k����������/�tc~N���t������1fb�����K>dU���h �!����ȡ>Muԓ�q�E�H��ĲB��Ta�-��L�S_7�	��mшt	G���J2ڸF����b|�Z��j/���0��	Da�u/��~E�^�.�'��]�K��SU`�Q�ho��mVb㱽�^\t�Ԙ�%������Xq�ؗ�3ݒ�V���8�e{�n1�����~��0��5�;��g�gSO=��]�n���U�'Hem�N4�D���L��w�����e�H� LMTib�#*Sq&�|����_Q$r_sv��&~��RfED�Y�Ʉߕ�4��K�ʽ�y�J�T�D&���0�R
��v�יACP���v$���)�h��Y���w���=L���2���iV�E�?D�&��J���������7&�=	h�|<�?�dQ���Ȋ&7�ӈt�(�է������)�������纫�/EP�����]!&J�D���su�O����4�aP@{�(��% B��f!��SY��@{�o�yn���n��c����2�fD=���^�+X��CG�ŴRd%��=��`KC�Al�b�O�B��~"�T|�)5��������^����D�G#�o6��d����yz�d�����=sUj�k��<�Tjz�~Fjn ��A�#����]#E1�1�ck0��/=�IP(�ml/D��i�X� �ɥ�$�l���.v�<�42�g��uC ��;��N��=���0��h�"R��Px�BR���Z5�05�{��/F���g��0B ��b��x^z����?_)c�bE"�Pd�'c{�(���A�)����/�DY�u�����a�"���f\�+o���G��G�Kx�J��{�5ٚp��?%u�\z�-+d��_�{�Q�W���'�ȭk��㖣E� ��g�҃��	�M��)�\H�}1V��}�����b�i#�?x��	Jٶ��+!�,�5�Lcb�g�����|�$�?�/v�x8){���Z��l�.A0���ˬ�iV6�����Z��/%��^d5�=���U�uW���bZ�|ƍwJ0����W���� 5H{��b�,�_�
x�'{���{���B[����`#\e���84i����U�`��oO*�#f v�n٠%�4� !f8H��*:#�@��8��`��b�cb�k��P��3I *�/�ޚsOd	q�dr�y��f-�+5WV��P���x�n�Ò�u_�[��M��3��^YZ�!���-���*�Z�֣��i�6��Ff�F��( F���S���a�LՀM�-����7�)ɔ���dӸx�N�;D�.Fu�i5��)�^4c�1�`%�#�v�@��̊QsφD9	��DyDw�>	�Qb3g��K�B'��S�4��a���^G�;�����p<�h�h�Ѣz�+��qCf�h/m�Q�׉�sJ�F��� ��G��]$Fb��hU��*p�����~�����n� ��Z]����m�@�c�Y|����b��EL�1:h-�4�t�C#���Q��X��7��^�X-�?+3�
�Z�t��/h�QF��L�L��
\��*y�g��ĸ��OC�� ��R��.�s����^�ɾ��_\H_��n^N�_, ��A���i7�J��P���p�����D��D�� ��c�4OD1�:�t7sF#܋� '�����P�B�Ba5����S��E���sH��E4��Ǩ�bYؿ0��؞ʌql]�������o!����y�.Z�eJA!�S�F�꫇�( �8���f����b K|UO���\��;G2R2AfA1���s$G��_.�

��bQ\�~�5�p�,&�v���æH�������Κ�2e���ȋ�&�'�kU�����Z���D���IL���)X_�?HK���aN�Ŝ��Cb������DǢJDl�:*>H�At��#��|v�uG3�<����7�nb{GS���J��ĵ��۬�"�-b��m�D���Ɲ[V��)��X�0!^!sA�8I�۪�B�	L��
]�R{��bLfb���Ho��b *3�r������xåTV�o?P��l���+!���Pc�1�43�G<�ޢ�{�v0��ڷXb{~�+��ᰘ��ia��Y�݈�_E��C�"�q�B d%T���]�M�qL�?1Q��Ru��Ę�f�;���z���MO�g.,"�GoS����%C)Vԗ�i�U�'/�a���ex+�r&J�#}�b{����Uī�5���p�.3Γv̌-jm#���AΓΐm����/�^���ۛ@�1L���()���Q� ƏҬ�Gv��zJ4=���W���t"ȷ�G&�j������'x*��-D��s�ul�-�e�RzV>���A@�Y5�4�eA�Av�KG�����nK��[��l�L�EsY\Q�Oϗ��?�X"�(#�R�KD1�rY�V�Gc/���6cJE�[j�v�!�{�5z��=���5%[(t-6�`)#�5ڋM���4v�	�ͬ�d��Ę�b�e�>���_<-ʊg̤�ɼq��2F����ϕRq茔͎���$V�TѰ�z��K"��z	b�ĸ��ak��b�!�jNe��g���ͭ��;t��T~�,sLj��b7��SX�����U�c{Qp�o�Ш�ߥ��'Һ�_�K&��,���3��ch���T�9Z� ��3K2zY���B��٣���)���( �	n+�l�����E\C{�R���Ȋ)�D�'����({�|kQ�U��Xi�E�;�`�k%�ߵHQ�u+��ki��OS���a���XW��)#��FM8���A�w�@���� ���D��(�T�Dy��r+����b��n���>27�21Z:K�ݥ�y�I�������n�9�dc������A[ (h�uۤLE����9�)�7x��4��_RP/NlF(�b1��v����~ 7{&�gQ�D�l�"Q@�ә�3g�1�f��b�%%�%�E�޼�j�z�R@�Q!���$��!������*�%�P�l���j��"F�S-D髋/l[�j{4,@�?ɰ��L�6�Xb��o�,�.5����RF�Kz�.�!$���e�\�R�jI��\Gt��D	0Q�:�=�)�8��qCeb�� �7E3BJ�l@jc؂���v��KJ���dePCs�����PV���_|�<�}UK������Q�$�����8;�NW�|2��obh�?�))x5��/��M�h���p������^As�K;6.�`�''��N*>���m&eJ��+f�{��|x�i��
F��R(�3��,]�Ĉ�@�N@�	$�Q����D� ��%��(��5c��O�޲-d���#7ÅdZ�,�V}Ku�����~O������_��[�%��r_�,������#taA:]��(RS+����ZAFk�������p�����є9���A2ڛ�F���/�D����O1%�'��-U{Ki��h�%ג��H4�e��J�)Z�p�����tߧ��U����ƻn�Pݪ2��N������U���e��b*9XC{U�s�����#��Gl֜�S�ьY��9-h��1�׏���7R6(�Cv�� ������5vZ����ܴ�&M:I��r�VҢ)z���V���LFo35��/*��~*���y�7��r��^i�7�\\A�m����K(�n5?6�ʆ��Sx�ץ74���pI`�jRv��oP���B�����DՃ,��:��k&�"��߀�b�Å��?߈�Ϳ���x�ޯ�h�<2�MYw=JP��)��lj���lAR�ץ��u�Xjz|���R�!S��)8���9�G�cO"��^C{U�æ�?�����j	E>�-h�Ί�--�$��D.Y�7k	�u��%� ;[G{%����u�8�쀌�H���1����'�>|���hb�t�?,C`��u�H��n��]d�i�����&�\�mQ�Ί8,���tK3M6rg��f��l��q����]z�������hozF>e �ݹM���
o>[���λ��Ƈ�n�`���Ϊ�hY���I��K�SA�l�@a4e;�i�Hj�odr�KFC�6���+�W ����5�I~�%�})���;w��d�ُ+V�������q_p����%��fy�F+ʩ��s�#P�(p�n	��MP�?��#]jG�4J��y�'��~�U�K|�uw�d�:��;��x�ukiϐ�G
�_�n~���p�d>v֛���+K�IV�24��a��;T3q'mX�5��L7�Lӵgjh�q3hܨ#����eA�@{Qa��D�%��R�j��>�$[+Z�C Mn؈���[�}�5�7҈7̼%�[u�����BɄ� C|r���K�,)&H1sãr��A'�ł�^#Ż�,X��k��z:��ǩπ�q�W�T��M�̣Q���%���[(�件�Zמҕz��I��ȶM���_"�)3'��������l����=Nڻ퐡R����T�{[���@�h/ʙbaeȕ7Ұ.��U;сBVkVP�̟	���D+���3�b!'�m�ᬀ�{��Q����k~�qB�* �0V��6|❌��	� ����Rj��ް���P<ȺS�7�iU_Y
��I����}{)�o���U���S�oj�u�T�Tf���6KW��?�*����dj��7���o=��+�fk�B�F���������o���$:q\	����*-����i�����t���B�qR3r���h�A����V�2ܒ����uiz�fQ$�%8b��~Ţ��\|o�.q]d�+��8�M�a#%������2p09�=Y�J��?5=e��@:�{�X]iHz���(�����Fq��-)�V�Pg
���<��wp�G-��J�߽���r�KA�3��a�����k	��U���?.���2A���ް�G� U	P���#kj�����I�|^���em�A"���n7�v�L~W����R��@{��j��䀴BL��'L��H�~uy��ͪ��D�>0��b%���RP���AbB#�����xx�Z�ab�E��[�V���T]@�]��噘����q��3���3�E#��n�k/�|�I/H�n�!lanС�KKU�j�ˢ)_,���5�~��ɨb�UŞ�<G�{��wu9�}�w+�@XO��Ȓ1�p�_"s�J;�<��M<��J�sN~+����D��oJ�;& �\h�B�FKXkd�v!*�Wz�	ګZ�J�yh/;�;��4%������
��8��Ye�=b<͘5W+#��Ɂe��������Eו��јC�c���\s�ށER�ߩ�n!8�>O�vZ7`b������S	�A	l���R�-���#0L��H������qXs�n 2B���<���R޷^��?�'D��F����饗����y�O$���֫��	"cS7�5�~�w9<z�F����S�'WJ���^�l^�a3����jbƎ�>�5�WA�Ij�HHd�U����E����0�;`�Illn�T�	.�/�W���4�)K#I�s>ƠpF���� ��̭��Z�>��	g�(�OOI|��'B`�
�Y�utU}ߛ���;[�HB`Gf��a�CM*�����K&�2F4^�HG{�yb�)DF�!3+�̻�5�j�?�L�Έ�:�/����N���>�G��DZ�s�h0���T/yT{ᙔq�L��(����9�g�݌҄��Ҽx�]|	�5�kdr�9��ЊY�����6��'�Ɛˆ���v�&/8D�a,���t>5�q���6��gk��שZk�u7�f{�����y���*m�����b�\�i�YS/���9�`�I�̻���e=})/���!��K�� �E�I/<y���;Q>~�d�p�C�r�������&��Q����n��D(�O���Μ�Z' W����7Ȕ�G��b���i�u��7b��q&J9+���C�@)���}�m���� w+��v�j2�� �`���5[Z�8��f��ꥱO;���ܟ�Ϛ.Vć}S9�>�'[�����)TR@
�����o}M�=Uz^0�oGh|�v�E��lb籣
_բ#����Y�$��5ڋ�%�b���{cװ��L���H2d �%� ���D3d|F)��H�ٰ)F���\�o[^��`pA�CG�C駀j&���,R�"J��"h/$�¹Z���U�Ǝ(��w���b�m�2g[�ETE����|1�br�Rz"
���Xw�%�=��JN���4o�*[-�v�����R�X��-B].H�����O"ˠc)�PF;�+(ĺ؞ʗ�HG
Pb������S�*+V�%O����z��#���c�a��_�Z"P��J+�A�B�1��B���+�(�8�Q�R���{"�G*p�^�>]}��}`v�������S�h�6v0�8%�U�7�����7L�/o=^+��,o6ۙ�-Q;�)T5o7����>�8
k~u�V�v?�V��i?����.|��q�8]�IEQ�Jp��M�����-�D�:��I�������`����(�o��>]j��/@�S����>}�o�nz�ˈ1�Y?0�~/l�9�����f��c�؟q}";�k9_�f�|��װ�.�����L�E�O$�k/r�w<�"������$�[��F�ؘr�I{/�<�d�v��,/Y!Z�ݕ��(:t�^\�=X�Y��_C��ְ���\( �G����4/����\.��e�����Ֆ.��8�t
�~W���8֐0�?�pR_zZ��'re=G�I�h/�����Tկ@�^ㆠ.v �$:�X����i��f��8���h8H��
~����v��(˥�=!u8�I<�D�H��U˨���o,�u���I��H���MiO�L�Q��
�fQ���I�zK01� ~7
K�O����o`��5��Ţ�~Nƅ ��y ��)������K��#@��YM�SI7��B�{Ļ�"l�[ل�0J�[�� I!z#|��$���ӦO�����>�$�K��(�����iDk�O���Wҏ��a,�@��}�aO��0w�ך#�����D��E{YL�h�.���)�m�521�\���᫷�f���#"�Ac�e����S}�29�޷��u�(C�2�i�H$ r2�NI/EI�<w���8uuk(��l�_�s�EYQX���@����jؑ�����kh��(%��z�Ԡ�!��V�8WR�^A���>y���t��z���YO���T�=�K�C:$�rLJ�e�|�� t&��'���r�qSE5�_�XGdy�+�)$RBW�+��1���5Qtq��n��:S��^�c�b��ؠY]x���d��a�W,�[�� %ak���h��ﱓ-����tk8��������F���R���ąx&T,�?� 88n���3���[�΍J3F&Sm#��Y�4`j;>�&���ġ���i�h2�iAr��4�P���Slg"�;�hXlKL���^��[����������c���XA-u,V!���dg���(1	�@U`W�֓P�E�'�z���^�q�菁àa;ofm��2c��x�dqh�r��ŦG������^DC<�T�u1b�;���bTD;�0�6�~i؛�K�����f�_�:c���8���K�9
�֮ ں�2�Q�#~���?�ܲY�!fsṅ�x<�m�^��-޺[�0>�t6�>fn |�.ab�D��m	h/���-� <���`Q� 0,-Q}�[hVJ�Y�h"���N�/��:�X�׫ڶ����4���`	����R��_�A��Z�n�eA{���9�n���<ـ���
����\�ld�i[>�?:{�I��b|�e��ޒ� ��iKe� _��0z)�'k/'y BJ��R�]X���Z,J�CF�Av$�8�՗/`E�G� El��I�?J�c����kl�<��G2A^2��r�-X%� %ڋ/&~�T��Y��G"�[]�U��6�YZ�?sFp�Dr_�[�`���lfV���/���n�/���#O ���h}G�T�V�kWhK��d��̙M���h+�z"7/�Wo����l�".K����=�4b�&���`c�8h�� �������7�qQ[C.~��uN�9����rP0�5w�#:hL��P) U�edb؀��y�>����|�*v-�(M@{���;�e���H���t��
;�If�t��#�V�`�m7ŋ�e�/���+6Q~F:��n
2!{+�!�LX�?��CVx�4��	�IѠ����um�������Y�x�f*�ʤ��t�5�߹��Ȅr%�=~��:M�x��]5��2 �^�g;�;� ̊�)l��Kt ��p�N
m�(N_�i��TUUQC%;>��a.ߪ�!Q[:��\D�ۧM�e=�ۻ��B,�3Ρ���4���i�ІhvQI��g3���69�Dol��&ې�F��Qh�z���O�ڒɁ����)��)\RB�!�w�]�]VFM�x�|sfu3�
ƐYJ �8ī�ָW ��� qDt�����U���d����u�{����FR�u$e�Tj��X5�)͞F��^��
5��lK���4���B^E�n��+��-o�I>�V���ʠ�c���G�A�g�����[���*�࠴�<�Dr�|������U�]a'2c�+M�_q-��Ss�UR��0�$o������z�vn])��M:x�hż���|�r�M�V��|�����)qx��5�}<�'��p������[Ѳo���Л�"�BA?m]����m�Sqe��6���xZ�K�7���_1�Ɂm���������%&��7��h��O��+o"��/�#�eM�o�B �5+(��MJ��}맷�Y�P䟳��?k��D��4�J����*(H+���'�{���T�eu�b���i�sΛ����+������A���Q<�����\����7�u~zc�<,�f�k�U��v2\�����kWhA�Xw����̪�?��[�;P۹{@���<�����tu���\�%��'��_����M���=9�!#L�Ŧh�����=۩�[Kӏ�pZ�L�H�|�FS&�"/"tEG*��)��j6]��]mlSe~����ʺ�cC ��}d�2�	"1$",$��E��	�hX�%� �?�EuL�&#sf�}�)h"$�#�97�n�-�]��޶�s��ֵ��x����=�=����9��D5��U�й�F��惰s�j>��r�3-�%e�N߮m�DXT�[ޞ*����1̴.���W �R�>���<��1�3���I6s=k"q��;H
��ywV���I�`*�d�L��+�g�6kBd.�l���7(yt+<{_C��S���ܫ�^��g���a�� 5�	j����N�ܛI�MgGϻ�[�߆����S���=�e�v��!�č�ptO����
��	�2�H��Z��~�p=?-I3HO��L E�c\!�m��h��/�n��Ȃ�q"e���l"�ڑ7�C1��jk�w��Warb���m�#�5���*�-�S��
�����+a�u����F��^ý�����S��l<�JKM�2^�U��IZ�j7�>2�7 #E?^B`Wb�Lt���� �$�����Km��EJ#�`p/��밷�O{x$�ݚ!P�n�-��`:�bf���_�[��"9�W�����]p:��e0�F��~!%��2Q)"���8���H�y!�Tp�����l6���Wj*u�]�dr3���8�W�Q^R���.��X߄��=��w>��� �~����6��D8z�d���{��аI
�3���n�#�d%V�B��$�tm64��Z��О�j!��-��������0�/��u�t��yT��$��b�V�!\~��B5�ll�cO�6��%�89�B�C����O�k�r
��'jT�l��o�Ů�\P���I���O��Q���?��G0�R8bF����a;| �������^�!���OVF}�#�3]_�r�u�͐�Ԧ0=2%npae�a����;ڸ�	���$�ىt����x~�š�P���mQ��"'� Wx�P��#�?6';O&�<-��z���EH�l��h8�J�*p��,B�7u9��X]�����s�8��3W�!����A��X��UB^�h�mu����}�a��s���9��6��:i�����&#%�o��l��n��\��X*c!�� {�~�Tw{���h4�2�sW̓��:W�[��"&�ي�/7�z�.L+I��KlN8C79v�S�[���:�ǑRb�=�����O���˅i��$V}�um��̰�(���,�\�*�[�h��Q�����(����Nz�Ø���8j���l.b�C�zE@��gޱ�� �Uŕx\��    IEND�B`�PK   ۍ�X���]  [  /   images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.png���S��i���S��>�����TJA� )��:��8I)�����Ox?�������~gؙ�$���@ �����#_>z' �1���<��K������������1I�n�g����q�~�����r��q�?�g�����VS1*8($Me�^]9�{ؐ���D7-;��ݣp����ԸT%�Q���%�B�ބqT��|>Z::o��x�A�4�3:߸�(ep�t����� ô�r���7�][7��G�ч���e��Ӭ��P����?�����dޏ�+3� ��O�W���U�����{���R0��Y��,��.����/ES�X��㺐��7���ZO���qlll_I�
XZY�ɩ�������/�?�?Dof 1�͏��>5U6w8��&(�l(�K��*�iyH��MU29��=�,���N�z|��;"��sQ�\BJ�<P�����kt�S"�*��ǘN�F,#�O}�T
kO��0?��s\�#������k(��u�д�F���]:���	׹b�w�)�5��b�r���D6x���NT�n�O��r�f��a���������JR�1m����СUPJ��1�6_��]���~Z���.����B2��Ŗ�
�S���Pp$q��%�O�k��[�ph%T�v<=9M#*����[2��}qA����h�!�0TT@���IC}o����	��� \Wv��v�霾�n��G����H���ե�ہ,2�D̍�Mhq�p�A�c�.P�~�ϛ�S	��E�F�,��J�:��@�EA�=��u@&�I�5���o�sg���J	���q`\y�#t+K��7��&8&�s8��$��ag�bY����L�:)p������m��9QG n>wU��	1cYNoqc�������'9����H�o�����(�:��_y��YS'��K��($H�XJ���Ox��\0Kr�DF�>J����z�?�7E�:�0������If��'S�6����Z��j�)��qZ(�>Tѻbz�_�J�K��sX��7vF�T��:P1������vf�C�a��+��,dK)�#���@�dy�\�ͫ2��zKB���\�,����2r�<�_u��^�U*�!��6ut-w5����e	L��)i�KG��I�L�r�S���`8?E� xaaV]����0���k�\&W������s�ؽ�*�-Y��U�=Z�����[��}�xOy����:/�P���r��s��+�w��׸�b�bm�F°�(�hj�l>b�S5��)���3��Oo��/?�?]e��F�_4T�R�0�}�u���{���iѱ�2=��CS���rLm�w��TA W��5^3�>����w���bܪ����%y"Mj\�2Zim������_�$�p������~�����~�:�������׉����w3(M;�ᬣ�L�GBҗVp�i�>�V�\.���e�êJ�/-{g�>8Z�w��E��O����ȴ��N$
��b��~���z����>P��לq�И*��L���ka��BƷ�'���̰1�W�)�у��#�|~B5w�5lX� �2�߬Bo8�s���h�I���ٳ�Dՙ#��?���:�Қ��+&�6y���hk�[�f�m�b��=f�� {�q� &�
ⱊ%�Ɋ��s���3���ט#�HA,��Ӛ���"�~�8�����#���q͞2Oz�Jg��`�"��*|\R���|dÙX�z���Q�Q6|��6��𱹻�����=�baf������������w�� Ip�8WB8���9��Th��ې�<*Z��/��' ɶ��7����d��� S�//Q��O��e�O���ā>y9+UJ!E�qg��:u�����5��{�������=Ҭ�Sd�l}*V���݄����aQ\���P��jO�+���3BѰ��:Y@����a�4c���ys�x���e���{ⲳ��n�mg�n#H�c��A��`�^X+����7KTVV���(O���熇�;�6^EB�1Gtaq�0J��m/�74+���%qF�6
�>Y,���ϟS���b P��O��D���H�;/ܗ766�m�p�L�a:�u/:*,$�%#���De����L9�a�M�ۓ������DTr���������z~>�s��͘.�[L�����͏�#�	nb�,i�3���7j����j.��v���5���WB�@��f�,��,rc!�?��αuZ�w]^9F5hC�444Έ���5���32��8Y�����S�l��[Q�d�ǽ������%� ��N������s��	�����21��33��#gg�CD^|�y&ʛ��E�:�e�����T��8;�K�;I3�IF�d�-gE�ao����z
a;}{rrrXUU�ܦ(��XFN��<=\ٙ�+�\��q���pR�{#&&��������&�M��� U�lv��όD"�!� �z@A�N��Y�j���_��^yz�>I:5�3�'[1b	�3fiJ��Wb1|�J=���gs|���"VK��II�p����w`[�ۍ"n�a�'�^s6����+�-rF��H��{���u:��d?�`6�l���$��`�O-5ޣ�w�LyÚ�t�e���ί_�����0?d� �n?ɦM�;~�}�T���-.����2'�z�Z��zS����%I#Z4[)���AR��-�j���z�/x^P�|�IR�Zg�5�ҏ��S�w�����Ӻ1@�V���D�JulM�z���>2Oo%LX+�IkЏ.��,��v[��0]vv�z�{$���P��_
�j�Z ��e��D���#�ͥj�oj�z/����6�$��n��܍p��4�D:g��'/�Ϙ��h�����f��[�We�\������N�+a�^�PӸBbXE ,D��*UPV�D} ���L2e���|�L�5:�Zjim��S��F�,F�E��w�B���0�ߨ����6�K���MS��:� �5�A�__�U!H�d��q�����1�M:��b]I�svVs����2}��a�7
;��y?�7�����n���Z/�Ifz��݁��/�*,5L��@n՛�"rT�[%��Q��}MpRG�����Qj�=1�=����'!��Zm��5���������!��U�>�#�5ߥ�(3}O��[�t80� a��P������-��Pd�����Q/��>O�\V�~��v���奦�W-u��5b��Z����1�i2�s�/_�P�����1	G��ks�"r��7�%s�jYL����_K�C��ɟk:l�����Ù��sP{����B��	xkJ{E�Vn�ί�_�4Q�/���/�uY���c�����cZa,ǅY�-��W&��]����*�n��Q})뵠�-+	���ڠ� �"SS���	+�"o�o��{G�ɛ���2*+�d릑�4�Y�ɍj����?KO`�Y�
���p�I���@��߄�gb����9|��wSp�?<��=�}�:��d��S9Փh±�Y�f�2S��ͧ��0�2�ܚN~�|W�I�2��b�PU�5�~��bm�F?�	-�V�zY��.\��U�S��veZ>��L�k�����������is��^��.���yz��t圕\�H0�3A,z�:~�Z�4�5*��Z��¥�������(;c�9�V&��"�Aq�TΠ�?��,e	��i���c�-��¹��*�x!F��Y\K��1�N�!���<�ۨ፩�6��4��'����K]Q>�<熉w��V=}��O<5��.ˈ}�}���y����b���Љꉌ�rdZ��.K�4�w[񧾿vf���pq�]@�e�me���3��޲G�zCBc��6�J=�|a3Ύ��$-��`9�w	��uT�0�����QaNMm0�H�5�[��DD'��s�!�����j0�6�ͫW;��YՋ��ͳ�ɂ
���a�7r���n~:Qفs�YU@�]�������#�o�$��/�Z3by.��R*��w־s����&QU���p8<
�S]GW��7j�Miˏ�-�/�:��?��Y&���*�R�̤�v?=;��В��	�JHHX�*ڍ5*�,j-��� n7������1��l&ۿD����Y�M����F�a�L�_��=$�K�b��Չ�}�n�z���O��E�@][��)�>�J����<;;$e���3.#���Al��ǿ�0���J�;$���:j%��'5h-�v ����<0	�4z>��e�r�A)]m�k4���[p�~{}Z |'>���#L�jll���W���%73�3����L�ޫ{YJ6~u��0�L�yq�(�,���r~�|4������Pͧ!�/��#�$XC�j
����o��(A��n`�ʳ��*
���&�?���Gs4]o�t9�	��zyOH�ˋ=��×j=��Bv���&��5�߭?�:	�� �� ���k���i�L�E}Vn�Y����ϗ?��'�Vo����{X"���BM�c4��(��L鐳�@����u1#>ǧ�Lm(�a)�RXۆ4�/�~S)�
Q��	@ӱK�ISe0�pj�?��;���fS}(�p�?����O��Nl꺲�ɟ�U���֮��6C���3�p�v�i��8�����p��)k˾�Iqc���O�	R�-�dy��k���!���T�tI1�LG�*�w��)z�]y
v�\s2<*��bA�IC�.Đ�����	n�!�wd{=����ϰt�E?�<R�w�_����pE�Oa�T� ��6]$r���^������)�~e:Y�&_� ϏH�,U:��`��@-�
���Fӭ�M*m�Z�X�Ž�I�4�C���b�P�AR����.�=����5��I� zÏ�=�"�	WNt�5�z�L$��Wn@�Ḽ��K�+]�_�"Ti�_-h2�
?��(�K��0�JG׮`�H�r����bGu�#�J�TJ|Ww��8\Wj9ͨ�~,I�b
c���M�Ƒýaxh$(�6ģ�|?"�l#ļ^�w�\CڞGpV^��X�~ۯ�	��.�);v��ZZ��(��ZH}O�y��[K��>S�垎%U�!t�,�PRjg�����#�pn3����\זM�H�"w�?��&nqt8��p��)��W���L�p���up-������t��	�ęշ���$�gP;i��C��u��w�OKn�S�W:k���~�4?#S-8<2 �֟\����Ӭ��=�D�>L�W��h�����@1�PK   ۍ�X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ۍ�X�Ч٦  �  /   images/e9f21cd1-5fad-45ac-b046-5921bcfe2a6c.png�WgP����Eo�*HSzI��P�w�׀�"����
R�P�HG:B ��4�E:/��b��;ߟ��qg�3��ٝs���;�s��Mt�h8i�������̮��Z ���xD��5 ��ldd�=�V�>o�k#(T�:�<�a(�%ă�DJz�"�\�<$C<�T8��h�������~��l����q,�Mn��XL6�\lq��'P���(,ql�Sp�R�ʊ�T%�:>��X����c�V7R����(Hr�?{��ln��`)f�C�`1��c̺�a��/y�Eb�R^�F*�d)k����6�ѥ�׃=ڟÂ�O5�G����Îִ���@ȉ�AҟߖNNE�!��WWV��YA��li��o�r9A�ഝP[���o� 2o�`�5� .-�,�(���m��$11qᲖو*�e�&1�Uw��a��22�j����B�-��u*��o{k�� ��F���c=�J�nŪΗ	��A���ԍ3#.��'`��`?)Su����$HK��6ཡ�<t��ֻ�`�J1���Ђ�����⨲�J`o��ۆ_�׏Гէd3���|��#�G�����<��8���R �#(���pvVO:v�R��`0�0��ʚ����o�Щ������B�*��͹T�э-Ty?4�jJ�ʏ�0��1���#��G\���>e�c����i��^_�,ݻ��	d�ฒw��I������+D }p%�&��
I_O~]d�x�h��
"w�n����������QQ��P����'�7D�d�L�| �7�ږ���g([��mof��#��CǺuI#� ӌc��"����x��0B���,ѻ��F1�%����y^А|5�4�{*�FON>ty`�v�~|��Q/u�$��\G�-9�1���6c�rK�Ϡ�w��z/�f@��\�(\��Y�	�F/�L�Y�\�'g9�żpI�)%������b#O}��[׹&���}!�6)��rqq����E��S�}Y&�\�GVL%n7����Qݫ�o2Vs�B�3�yԚ�k)w��J����fF��zNM���a�䷃z;�[f��A�u��i�&Hrb1����"��w��F ��}q�?��C&�L�j{A�K鹖����/G�c��ݍ�1�2�z�g��i�aa�c��A1�vޥ|�_��	j����Ǝ��[EW�T����|�Q���[��=�x��� /ÛJ=�a���ՙ�ouc��p�;d��-F���;O�S�Z��{�x���}�zOBa�����G��GwP0����7Ss��Rch��M�!�)�RP��7ZR,� ��OS�Z�]��r2n�f���tS���{�ۘ��	b�ڡ�]s����|)�fok寜�`<�}�upB+v�C�P��$��]N��V��!�%���:�i���+�>����:,��$��Ot[�)�hMy�ͱ���9��B/x|��j�:(m�꺂��]��8-0!˥ʂ%�����Z���E�� �B�U�yF�ڷY2�񛣣��㦿L�H7Ű�߿P���^��b����j�׵766��׼_XA��]^�մmmF��(E�XN4d�����\!o�}@۫J�m"/z��}	6UUU%�@�⿢��ٵ��;��X�.���L1v+���H�tO�`l����4��^�D�s����B���*b��++&s�ͼ&ad=*�\��Mֺ����{ԴF��f1K�=4�'?fgK����3J2x�6d�r4HK��"�%2�X��t�dR�ٵ`�Xr���}}����#9��O�\7a�\�o�'7ܺ��.�jad o9PA5�77j��I�o}<�tx#�`��Y.����Q=Ӝ��L��JP;���}�[��>����m�^g ��<��+0[yr���ӭ��M�	����v0T��3������/��]���>�î��
����T��WiU�����.������.�g �l�ss����y���*k�E-'\��Xm?b��������(��Qx�v�`x�č;��֮�������l��9K��2S:�[�`�񣣣���E_߽��*ܕ�w=�)b�L�(Y�H�\:qONMMM����CM��9%�2����?^"�@��1�Ki'gf�<m�3i\�q�b�_�K�xy��ڛ��H�:�1[/�P�\�p�g�,r�+��$m6��1�OV�/�ј;���q�j�c��_�1�*�1(�����&Ƚ,�"�^��}�Z'"�'��籵�n��2��G�|~⬋F!�c�@
��B,I:�]I�f�JlL!���ȬU�!���\Y���v5o����hx�w��??Xo�B�����09��&���:a�<�(��H�4���b@)oiYn���/C%F�NN��W��x����,�\wi_��X,AG``�����-�+�mO�|�����i�L�=���LBB���H�a��/V���#���c��.�S��9v�j	�V����������'��T�9��Vb_����6z�('���A�D������F����e�,8���!&_�^�(���I�0`5uW`x>w��`�D�1�u?�G�TB	e����6�d��l!2X�Ͱ>�v��4P �H�W�RQg�����7z�v�	#�_�(�dM�-�č����qy�]Sy�A�,�P������V6\�k���Aw��|��}X:��T4+l�FK+�����)�ȡ2c��v&f�{�8�H�f�h���t'�C�����:���ҬKRo���E����'����{{8�F}f�z����bOH��l7�X���z����<K@�t�O�o�3x����%?�yY�d�H_��8>8��t��5��V��K��|?��k;���c�ڇ��vUg�ǹmQ�:/��'a�?���f�|/���d�:yPw�=��������	|�j��~)�H��e��/�Z����X���X�C.�Lm��|����N7M��5⁌-��eVs)>?����箷��O�aW�C�<j�ڟ�sx}!�l4�YW�8��j;j�>3Ӭ��"�v��8��� ���H����hO�z6�U�OB0 ��d��d:�	��Ŷ.��8>8D\E���/���y�����������W)̴�V�KKC����p�5��?�f�h@:���Ԩ����\#B�V��q�A�TV&d@�!�\o���2�$,����:�+2s~����뙯?*d��&Z�0�PK   }��X��/H
  V�     jsons/user_defined.json��n��_� ��P3}�O�ĉ/H^���X�i�f�<�1?P^&ϔ^:�RZن�kH6����W%v��S��"��g�<�-�2�r�����ɨ��:��Lf�i:�?�����3޼�����Y�{1�{OGq\C���]=��ʬ�=�.�<,�l��#��'�ْ�%9[ET��Xf�6J���e?�yǣ�颓�ϿExK&%M���l�'���DA������bT=�J���_�·��ř�x\����̀q*��|��м��@[��BaqTf�����z�N�����kԓQ�ѧ�3xF+8���[lr�F��*��������x��ܼ̇���u���v}֥O�������ٰ5 ��[���?yt��ek��.#�^���}��7;�E���_n1�K����y���u~Y��鐗K���yS����y���unO��٪�:��rK�����y;_� K7p�Ϯ�O�G�Bx���Y�)`��T��w������=<C�.�	�Z~��;4������C�.�	�Z~_���]~��3��5e��&�k�}�m��l�ݵ���<l�M�	�Z~߬ҙ7�]��;�;��;���i��Enker#��7`�o�5��E!�a4���3<5�/�x:Z���:s�բv<���rӟ͚G�G��Z6��<]�v��ϫ���b��"_�&�p��ύ��y�y���v[L_͊���8��_�����(�բ����BI2{"��$8_M)����-��q�*W�W����ҹ���PP/��3�<�-��>�O��b������ޣ*�i�{W����l�Y�+���6��"!sAD�-S��	:_�߷
זj�C!� �J⠐'*�Hs�^{�G.�:÷U�j����P�3!~쁠�lt����	��Գ)����|�ʜCPGaW���i���.����8���x�~!�H�9?�n�,U�2�e��k{y��}B.��x&_ƳѴ��J��=��{&�h���x%�V����@J)/�H:���#�!�p}ʽ��tZW�v������yÝ��C�a%QE�MF���X�]�r���<M��Hgq��]�.�d�U{ πy�����0Ɍ��glX��d�1*v|�VսfL�>��-0�Rd��U�y���ݵ8��4��K�.��Da�Q��3�1�s.�|1�>�M�FO�&�4�)Y�M�D�TH��#�	<�\%&[N8�d��8�"	�jc�-,h$��~PҲ+��Ĉ*>A�a�Q��r��X2�:"iH��]��n�su'҂�%Z�I�,�M$�Gx*4'sta_Ҙg&��HQ��zQ�V�T&�t�I�j���4T�,k�|���"N;E�HZZ�-��9s��:�!iH��EH;ɓ�dZߜ^8�����犐YP���l�R�,EJmT{O%x-���-`� AE�k���b3_��6�������ԏ�/��_��b����4s�n4[�=�֬�&�K�,��/�uewOn ]�s�6��n���U&��?|3P[�L��y}��b��*�KJ8tv���s���q�����t�w��_�i���<t&����/�<���~��|�5��%Ο���54�������f�o!��,6{�lv����|�&�}RW;$ԁ�+�5G�"��R&4+	���^�P�.������������������_�p^?��y�1/��s/�^̽�� {0�z�8}�;��*�Ms����\yD�*��K`[��%�+�<�6�G��^}1 ��΀:�4D�dIcD�y�3m�MΪ�ՓW��2���@�N�'�Hb�D�3�q�]n��J+T7���n���F�6�nO�EZg��o��m.@�?��˒����B�~{.�ݹ���##�Af�J�`���n]qPa��6���	VDs#)�d�O�!��%�6	w\�{�¨/��n�?����o����r�\ �r�\ �r�\ ߖ��,�A� �M� �!�w����sy��,�A��<�A� �w���"�\���Ep�::::::::::::��'�q��{��F.���@.���@.���@.���@.�������q�gnp�f�O�^~��	���u�����T� i�%؂*��R$�@�u�&�/���0���;�vI����EP���X�	$dN�b�,u\� �|��]�A�m��A��6DH6�n�7�^��S��=@ Gwt�Q{on�����f|��6[mB�Ҋ��,�Wk��>!O�(��/���r��k������!���!G�����8��q,BQ�!�eUJ�qE\W�qE\W�qE\�{�5�~��jk<��w��!�PaR�ݝV�4��b�?�)u��!x+%�i��h����/��Q������[�z4�}d�ؐ��4Fbu�D� P�\�(0���Q2���]D'�%�,X$*�I��h]&�(�e��swb��6�$f�޲�J琵��ZR�RX!$�}+5?�6q�u�Dg�`0��:ʓϹx��$��"�����*N�n��uqZ��uZ/��EҸH/@.��x +H� ��Ŀ)�����#���?PK
   }��XB�*h  ��                  cirkitFile.jsonPK
   �{�X�����   �!  /             Wh  images/00133a18-aa29-496d-ad09-d18fc42e20cb.pngPK
   ۍ�X��`H�  /  /             p�  images/0b5b01e6-dad2-4c75-9695-e3d6481bcc1b.pngPK
   ۍ�XK�`��  � /             ��  images/1a17dab1-c3c5-4679-bc59-2ce04d496e8a.pngPK
   *��X�����   �!  /             �s images/4b131f3d-bb43-41b7-a007-3fb3641e8d39.pngPK
   ۍ�XS�ѝ�  ��  /             �� images/642b7e82-22f3-4f40-989c-bd067878f1b6.pngPK
   ۍ�X~��k�6 4 /              7 images/663b53f5-e86a-4272-a51e-f5b809259b46.pngPK
   ۍ�X��L˪ x� /             �m images/68064abf-29c0-456b-9754-5c6c0ecaa6a0.pngPK
   *��Xj���(  *  /              images/6c8b06c1-8935-4e1c-b7d7-4989f9141afd.pngPK
   ۍ�X����O  J  /             -B images/76768ab9-a537-485b-9af2-6ea55daf4943.pngPK
   ۍ�Xd��  �   /             �Z images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   ۍ�X�1.:�  )  /             �z images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   ۍ�X}�Ί  Q  /             �� images/a41c66fb-6d0b-4037-a131-23cbdfceef6f.pngPK
   ۍ�X	��#u } /             a� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ۍ�X+L$��� �� /             �	 images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
   �{�Xj���(  *  /             �� images/b092be47-6ed8-47c8-af5c-3a16748d9859.pngPK
   ۍ�XᎩ���  � /              images/b3182cb6-763b-4979-9bf3-a9ce9c9d7585.pngPK
   ۍ�X#�@�9� �( /             H� images/bb1d7dd6-69b0-4e8d-a72d-bbaa9fc3070c.pngPK
   ۍ�X����<  �  /             �� images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
   ۍ�X�ĩ�xa  na  /             W images/c9c0af01-d4ea-463a-b9af-0ddeafc58269.pngPK
   ۍ�X���]  [  /             f images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.pngPK
   ۍ�X�GDU7� �� /             n{ images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ۍ�X�Ч٦  �  /             �^ images/e9f21cd1-5fad-45ac-b046-5921bcfe2a6c.pngPK
   }��X��/H
  V�               �k jsons/user_defined.jsonPK      �  bv   