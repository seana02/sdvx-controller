PK   }��X�,�KƘ  j�	    cirkitFile.json�۲帑$�/9��nA��y����m㵧lJ�e��ִ����wVW�Z�8�[:9f�]|9�` ��ç���_^揟֗_?���|�����������_���?}���_^~����_���?�����o���j�O�L˘�%u�د��|7�hgg�ά.G��bx�/�ß�"���S;�{% A(���	/�k�~����|����ǟ�O?����_Ed��)�yd�+��!�{E�ܝ�� �~����D�\�^xGd��B:!'#���*��s`* #P�L��K'�4bK	�^�@΁��
��[��
�[ ��R�P\�i��4q�1(��XY�V��4��B�@�%99Da!˓v f�褉߫5�=_��޽^�,[�͑�:�5$��J�ܽ�^Q/b�9�8�Jsa
���y���Q
Qt����[�g���%��g��w��Q�`ϵ�xi�(U@F�5�	su�����w���ξ*37��4Oqr��z�z$~Х��^��89Da�K������P�#q�$ݼ2p���uR&�t��@Þ>��%H�`��K���H����6R�o
�X����4�	��3�>L���#2�!�]j�&�p!'篇2	��_��P�L��,���D�U%M�C��1)��O�.\��J8�]�V�89Da!+������.	3zDq�#=R2x=�j�O���GȠ ���Ϻ4m���
	� �Y���99Da!�0C�}��YHs�)|�'b��B~"%��/�|�C�m1Da!��Cr'/�(,�b��Bz���<�!
y�C��)�(,�Sa_�<v�!
y�C��y1���d�j�l����9�����Y��n�������Å� )��z� �k�A��������-)��{2R��7d�o��2R��jx)��zta�"D��j+��	�!c�j��C�;}�6%�"���d;�VBA��;��B������]�@�b�5Ua/��Q�ǡh�9-�A/B�,�!�
��DO���u�E��١Y���1o�X1��i��|��i�:EdK��jy�E�3��;�"NO0a �]%8U�U�r�*����FY���ye4�����!_��i�|/���y�:���r�h�zNO��)rZ&�^�<�8/����"���b�h���7&����ۆ�u��&e!�����.�{���υ�" i�N_����Y�/�b��Zd���H���4�֎z[eV�����_��� ����zd4|���!?2C|.H���N��s��K{<}�
`>�Q�&D�	D'=���,#JO "�"��⩨�iSTx2���B�Y���o'epU\��5�&�Wu��c^���_U�!_���u�(�Ͼ*��s+٣u�Z����I���w2ы�-�; ��*�|;���e!��ճw����x���4�� ��6���+�UQ6z���(e!_���Q��(e!_���Ab��n��|Z\�}]���Y}����̐�d��f��8��|]�!\�u�.�9H.�A�{q�����u� )�e]7�A�pY�r�"\�u���u� )�e]7�A�p�g�ԧ9���iO]N�\Ћ8=xE������<�_B�,�����6�B�
�Q�Us��8ݏD��Ӄ �"�K��^V��,Nk�P)Ow�Ћ��:b{Y�楲��]��!_v���(y࿪fEY��U5+�B���QQ�[]��>ݯC/B�n�!�e�&�B��<��!��-Q��}U+��yq�>=�F/B��WMh�M�C~U�nH���uZ�"��F8=A�lF^h�!_v���e!_7�*	Q��!��ו��Eȗ��JB��|ٹ*DW�F�U��B�n\�ߡ,��U�ʂ��O���:������_�_~{�֭�r�&�a21��i6�[�m����o�I7W�
���y��{*���q^5�o(/B��W��L��P��RB�{d�a��j��%^�}Nf�q�y�~�!<����jA�lK���HF����@�l�!�Q�d�?)ʂPF@�#����:6����]ձ�,���Wul(�Q��cCYȍ�U�Bq]
���5q�A)\}�������d��s\ve�j��Qٹgv�� ��s���kۋ*eBS��=_�L��U>p��;�$�I���;��G��Tv�ˮd?\�:�vTv�ˮ�)\�W;*;�eg_z�v=W;*;�eg_2W��Վ��q�ٗ����Վ��q���r䴞쉸���^oO֏��ƈ��~�>���82��v���%[���Kܡ��
�幃��E�)�����Kv*\~_w��G6+��$ۋ��qO�B��'�F�#ۥ����Q�';�����%{&.��-$�~d�������W��G�N\~�UFs+��'{/��mD;���s��s�'��l�?� �^�u���߶#�G�n\~��oO��|	s˯�P�'[7.���RA��d�������W;������#�_}V���<q�=FE�|��pG�^��ۈ���������	�"[��Ϲ���lݸ��7�������#����f&_Aj�����xx���+����;�'Z��t#[�@�n\~���~�Q#�~��@��z�'����5�E�n�����9�幃��Ev~�ߒ_/��q��}!������#���c]��M�$�&��lݸ��^��K�n\~h����d�������W_1��Z@�n\~�_m�M�(}�)��_$:++�<G�<wpyB������s��%;?.���Y?����sd~{�"f��N2�_c�F�n�l�"ٺ=�-VR'ν���Y~����sd~{[)�~d��������Vd��֍�ϑ��ݰ������#��;iq���ދ�ϑ��]�����͸�����>�x�����~�aP�~d�����!T������*�^�}�������c��`7� ����?:����sd~{�=�~d��������d�����ϑ��}������#��;2r�Kd�������^�d�����ϑ��]0Ϸ7�=��Q��Z���q��V�C��c['g����ch�>��p�����.�.��chGe���/�*��chGe�w�/�&��chGe�w�/�"��chGe�w�/���chGe�w�/���chGe�w�/���chGe�w�/���chGe�w�D�Y����_��,�Zp�Ut�l���Ƕdw�l���G�����`��m
T.�G��_�Hv)\~�9�(����3?��=��D�"[����g��w���G��d�w�D��엸�*�s6���i T.�傛{�H6]p�L�zɶ�˯��gE?���{�h���~ـGٜ'[7.���x���홟d����Q��GK�%���t	�~ـGяlݸ�*�s6�ɓ/�?*����=�$[7�y&z�d���W�ܳ���{��=a4��E�np�K��ދ˯�;gE?��z�'��Y:}��n��^ ٺq�5���Q�{�ދ˯�;gE?����h�ـGяl���*�k6�Q�cW�a�5a4����l���O6O\~�1�(����3?���ӗ���������Q{M�|��"*�{��5�${/��&z�d���W�����<q�U��l��T����F�^p�<��d���W�����{=�M_i�"���"?ٺq�����Q�c�\E�^p��<�~d���Wѡ����<q�Ut�l���Gv?\~*�(����_E��<�~d���Wѡ���~.��p�Ut�l���G�/\~G*%�e�4��H�r���_E��<�~d���O�;����O���I��^^E{M�ٽ)��)��)��	n_ـGяl���*�k6�Q�#�'.����x���˯��fE?�y��h�ـGi�C6O\~�5�(�����Q{ME?������-.�dV_@�83�-�4��v1��8��m,�����6��p��G�������X����chGe���/���chGe���/���p���6��ŢV�������XԆ��1�����X��Z�z8�vTvxK�bQ�]�Ў�oc	^,j����Q��m,�d�l,�6�h:K�\~m,�(����_�m"�(��-�_E�<�~d���Wч����jp�U4�l���G�\~� �(��-�_E'�<�~d���W�ʱ���zp�U�rl���G�\~��(;�d���Wы����p�U4Sl����>� ��YaE?����h�؀Gя�?��*�!6�Q�#�.��n�x����˯��aE?����hg؀Gя�?��*�6�Q�#�.��~�x�*�����G؀Gя�?��*�6�Q�#�.��~�x��eVd�7�k���G�\~�(����_EG�<�~d���W�����p�U��k���G�\~-��(����_EK�<J�3�p�U��k���G�\~=��(����_ES�<�~d���W�T����U�����5�Q�#�.���zx����˯��^E?����h�׀Gя�?��*��5�Q�#�.���zx�����˯��^E?����;j��ã�G�\~]��(����_E[�<�~d���Wї����us�����5�Q�#�.���tx����˯�/]E?�����K׀Gя�?��*��5�Q:n���_E_�<�~d���Wї����\�?��׏�����R��y٢qn�&nq4��73��s�aٖ+�dýlx����lx��eól� �6�i'�wN8�p�9��s¹焓�	g�N?'�^8��4�	�?��/�o1�q��_L�o�!-��c�Bw����W�4M�8��ٲ��5�)�֔��a�y\��_������֯���kW�`M�lW�\�4�eu��uh���O�ݺ$�5�7��r�[CX�u�Zo�����./��f��B~L��2��5uqs�_�_�����2-���lư���+��2}���D��x��������:�2��s_������j�!�9�<��^�wd�ů�`]��N�d�d}�6�jV��-�c�,�կ#��=�n����~�ʍs[���<A>�	[�Ik��'~��q�\_�f�S�l��r	v6��Ӷ���i��uh���wq^���H��n2y�:3Nۼ�˚�>\�:4��ׇ>�q��lc�o�L����q��S��uh���ϗh��*Sʺ�u5����}���ά��؏�u�ŵC�ϯ~~����k���R�y1�LR3�љn�cZ]Y7��kG�_\;2��ڑ���Ѝ}J��S*�җ`���o�}��1�4oW�~�[!�/R+d����S��/���Ȥ�O;���5na�W�4��ڡ������a�Bߗ ��ex��ɶ�G��!t�d��j���_�wd��}G�_d�}~-+�ds�6%3ô�����O���4��ڡ���?����JRF���H7�呉s2�T��4�yخ�wh�EN�?�vh��}湟KB4n�X�i(�KJ`J^�ء/����i���~qߑ��׾,[�G��q�%-�s��4�)��w%?�׫5~�&����^��4�|�~�}?߽���o�@���n�i#�v�yw�w��μ��Cl�p�]�bㅳ�b�/�{��xi�ο��åOn-k��R˂�%3x���a�n�[?]F}d���#�/.~~�s��<�b
�՗�}4Ӿ�ִ����G�d�ϯ~~����k�<:�q�+I����>y�}̖�s�l��;����d��������d�ɕDi�3&;�0�~�Kr�*˃��_;4��ڡ��v��h�Ɍ�?�)�J�8�h6�m�9��-_9Zd���E�_8Zd��NFCv�t�/�L(�R��u7�a�����Ch��N0�j'~�ꖸ�Ώ�<6n��E��]��]{��C�/\2���!�ϯ}K��,e��%Tv�,�E:;,��.�0^�wh���C�ϯ~�A�/ң4-��f������.e�m�(_����^� �/�d�Ez��H-����ukI?r.KS��8���llW���ϋ�W�4��~.4�������h������[h�������:h�p�]�il�p޽��?FO��q�>���}���N�;��N�;��N�;��N�;����Maܼ�����<w��J�SV������CYɇe��|��_������~~�O�����^��V��j�[s.6g+��*E��_�5 �ϯ~~�n�m��^~U��h�hƾ���ݼ�1�y������.d���C�/]�<l>FS�M��Ӹ��gW�MrÔ��;wu��8tA�_� �/,�8n�K�˚�t}.F>g�e���ש�����K�������k���ݘ�`y-�L�����ޤ-�ɏ}���!+4��t~~����m���!�g�C(��,f��d�4���K7��9��U��_����i����m�{�継1���Os��ۦ0]�@ï���׎������(�qC��eIEy�B�6�3aۆ���c���C�_,����%~.4�\�0����������͐J��[��M���
F���L����D
����lƒ�d��S��tU0
�*,�ð��)I�j�J�RR2���w���We������-�e)����&��XN�++��}�w�%����_����/�}|�?���Ӈ?���\�s6��^d���JY��/�lu9�u����ч��m˔҇?��7 ���$@������6^������Q��s��C��ro@���ŷy4�~�1zZ��JZƨ{�Gn)~E��hZ�0��v�\����_K�="v����k��Q�	#v_�]���Q~c4���;���<l2F�@��,�k�s��0C�+�T��Dg_7KwN�* �#ž�mG����d_we9��#-�u����!Q8u�4��qJ���}F�p�is��ŧ�؛rX�p�}C�/��u7��	ɾ��K�}=5�ܻ7$�
�=+�|Cb�qOʜi��&k����oV��;�Eȩ�$��w i:���i������v�2����e�ސ:ˊoH�m�����mG*���q�In��o��t���!�bi����u�݋�X�oH�zZ,��L��$��[JoHyf!�������i��+�������c�)֞��H���Y����C�6�i�*������o}�8���D��,���4N�}���YH��h�h�xG�g!�=�i�h�xG�Wa!��i�hq���q��3�Ɖ���!�q����YH{�l'�ރ�Ɖ�-�Hs�1L֬v�&�ٚ�c(�yH�u����@9��������,P2�ݵ�%dD�\W�`D�\W�`D��"9#�����>�1��>�1����+"�H^ԾߵB9��G�msg��('Z�v���(���"�-v����	�"�@('Z���PN���`\Ŝh!��d�j �-���Sd�	�����J	4���qO��,���(	8-�������hY�[5P�OggP('Z����('��uE���('Z���DB����0�i�x���,$���D�G	�8����ys���,���(:���[5E'�E��PN��@��ߐ�eN�5('ڦ
鏺"���K�,�ä��x_�r������_~�"-�GھJ���,���>8F�~A���G9u�}��j �G �PN�|�PB9��8	�+B9��q�=���5�B99V��VtY��r�� �@('Z>���ǻ��U�j �S���j �-��@('Z��PN�8T��hq�B�i�*@5ʉ��ª���o��6�%!uE #RW2�ݵ��dDB��&�,F�/Ȉ����H@H]Ȉ����H@H]Ȉ�{]�e�4D�6/l�"]��r�o/�mG9�"7P�r��n��ʉ��j �-~uE(�W�5w�$���B�H5��B)o[w�n;ʉ�YH�B�W����(�D��,$���D��@5ʉǁj �-��@(���_}�z���hq��d�j �-�{Zg!AuE('Z��P;��4�<�Yȉ�YH�]��@9}�`w�I���J���j�a�6�PW�r��q�E��PN�8���^�.;G��hq�����hq�+B71i�*@]ʉǁ�"�-��PN�=qަxd� ]�PN��PN�8�����@5ʩg�a�U1��H�<��j yN�����H�����X�?W��G��@5ʉǁ�"�-�]�PN��M��&-��PN�|�B9��U�j �-��PN�|�B�i�8P�r���j��_?�}�d>�?���׏?��~��?��)����+թpu*\m���թ���p}���W�����:��+C���kP���\�k�E�D]���QEW�N�kɃTt�Tt���T��EEפ��W��վ�*��*�jpu*\�KV�5���թp�/������\�
׽&X��8.�N��^۬����R�]l�mm5܌�a�t���:�>;��Ua��RD�1`Nǁ��u:l��mu\�[ƶ�
���_�2�ձb*l�w1t歎Sa�t����h���T�:���1:��2��-�\AǗ�g�C9Y��el)"��2���T�:��;W:���2�N����J�uN�زa����2���T�:���|:���2�N���N���:�L��;bK��t|�v:�LǗ�����˼�/Sa�t����h���T�:��;�*9X�9/;`ˆej��˂�/Sa��2ֲ��˂�/Sa�t����h�T�����R歎/�N�����uGl)"������T�:�{�mu|�
[��v��霗�e�2���eAǗ��uGl)k��/:�L���a���P�6��2��-c�F_5���a��RD��eQǗ��u:l��.:���2�N��ޣF%�Jo�)�J��ˢ�/�:��-��Q���3HG[_�����{�h���T�:�{'mu|�
[��v�E����/Sa�t��=�T��t|�
[��v�����y�
[��v�q����/Sa�t���t���e*l�۽眎�:�L���a�����V�ˇR�_����NǗ��u:l�^�:���2�N��ޓQG[_�����{K�h���T�:�{�Lm��/Sa�t��>u���e*l�۽g�ʹC��e*l]5[�;ӕY=*�ku��zT���X=*QW�G�W
Tnzԣu��Z�{T�rã�����ޫ�����D]5�V�^���G%�����*�@�&G=*QW�սWA*78�Q��jp��
*P��Q�J�U�ku�UP�ʍ�zT��\�{������f���:�K�m}��X��J�K�w�v3m�ej�c��^V��"蘯�n��:�K�m}��X��:�-e�꘰�n�r���W)�����n���y�c�T���^m�e�[;V�{Aǐ�v3EEбd*l�{�6�2�ձe��W� _V��=��e*l�{�6�2���el)�V�@L�DL�HL�L���i,S[_�¶��j,1Sa[�{AǗ�v3EE��e*l�{�6�2���e��WQt|Ym7ST_�¶��j,S[_v��2ou|Ym7ST_�����*�Y����T���^m�ej���T���^m�ej���T���^m�ej�T�X�{AǗ�v3EE��e*l�{�6�2���el)�VǗ�v3EE��e*l{��a�{5*l�{��"����ޫ�:�L�m}��X��:�L�m}��X�:����**��/��f�����T���^m�ej����R歎/��f�����T��^e�2�Uz�LǗ��^m�ej���T���^m�ej���T���^m�ej���T���^m�ej���T���^m�ej���T���^m�e����T���^m�ej���T��^��� ��VǗ����� ��VǗ�ex��n��Ľq���WQ��|(u�Pj���j��6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2;+��2���W`����2���WٰLmu|Y-ې�����v�g��%�f7�.�q��ޫ��4�սW�Q��V>`��D]5�V�^�|��Q��jp��
*P��Q�J�U�ku�UP��͎zT��\�{��
Tntԣu��Z�{T�r�������ޫ����D]5�V�^��ܨG%�����*�@��F=*QW�սW�^�p�v3Esx˥¶��j,S[%ۥ�j��6�2�ձ^*l�{�6�2�ձ_*l�{�6�2�ձ`*l�{�6�2�ձa*l�{�6�2�ձb*l�{�6�2�ձc*l�{�6�2�ձd*l�{�6�2�ձe*l�{�6�2Ot|�
��ޫ�Lmu|�
��ޫ�Lm���t|Ym7�X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��Xfe��/Sa[�{�����/Sa[�{�����/Sa[�{����R���/��f� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� �|�AǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��V�U2_V�ʹ����/Sa[�{�����/Sa[�{�����/Sa[�{�����/Sa[�{�����/Sa[�{���f��/Sa[�{�����/Sa{�{���VǗ����� ��VǗ����� ��VǗ����� ��V�͇�/��f� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� �쬤��T���^m�ej���T���^m�ej��� ��ǿ������^�H?/[4�m��-�f��f洹a�6,��b)(���)(��)(%QPz
J���YG�����8��q��L`Ǚ��3�g;�$v�Y�9�ؓb0g��Y����i0����n�f�:?�.t���r����4��h:g����h�4ZS�oG_�q��@(�\|�~�l4vX��k�d������d�=�˴�ЭK2nYC�"כi�K��ޭ!,�:�r˥�]^z�Ͱ���4��+�p\S�1��u����rY�����q���b��0�>���>w��r?_�]�\ �9��q���e5ːҜb{g�����s���n���M&N֗Yׯf����<v�2\�[.�vS����kW�������S��%۶v�i�K�7ח�^nm7�h�\����`��mkvs�@(�\�8�~���Eݡ�LަΌ�6/����\ �[.C��8�l�1�wz&�C���_��)�s�P8\nG�vm,6p�⺚���ľ��`g�u�k��ٺ�^�V�V�^�-�.����ˌ7����>�Օ`CtAP�uAP�uAP��Ѝ}J�,hS*�ۗ����o�}��1�4o��GP�L�>�DPnu�0���7Ώ�iLi�uv0�-�k��B��B��B��/a�Bߗش�%��d[��,$!t�d�X!��������ޓ�!�����e֕���6�~�c?��2 9&�r��r��r�K�u%/�Y�\���4�9�n*~"v6 �P�} �r��r?_�y����/�s
J�|LI;�%x���P���r?_�[]�e���V3αd�q.j�f3�����y�i�ޫ!(��@(]n7� ��};�v�B�ݵ�Pn7� ��=;l֑&/g���<c0��{���pf���3Ù��;�g��<c0�̙��;�K��Z�63�4��Kf�6g��ݒ�~BV'�^�^�V�9�e�C����Jʹo��5-k����R
ʭ.ʭ.ʭ.ÐG�c6nq%��]4y��ްo��2�	���R!(��Tʭ.)�!�0�mr%WܦŌ�N�xM���\�_�V�V�~�a��h�Ɍ�?�G�J=�h6�m�9�b4�]�~�A��u@P�]�4���B_��P����u�����;�
�K� �T ʽ�^��:?��D�}Og��<7tѮv,_ �{w��ܻk�V�-y?ز��U?��ݹ��u�ﺐ���V�V�6E�P�3�4-��f�����.e�n�ܣ8����
�a"(�Y�r�!(�	8�r�n���+粮���ġ�+fc��wl~^�rL���A�UB�}�!�[	���G��>B(��B���
g���`0������n�V	g���`0�|���p���Ù��; )s���ȸ���n6[I���Vrv�`�ws(�Ű�y�r�P�{��������y��0��G9mf�5n͹������!���!�V�V��6�m/�,�|�c4c_�h7�mLy^�����j"(��@(��s6�)����4n&�����0ek�������r����;�q�F���5u�l����mYg��u����#(�NA��e
�wc.��<��қ<�ޤ-�ɏ}�P_ ����"(��@(�;��Cܫ��L,+��z7�<�ns���x� �{/���{Q�^�i��D�m�{E���1���9��mS���.�yP�uAP�=:�r�!�1�c��,��#�B�u�3aۆ���cF�r���A�_��[u!�[uÐ�n��r�⚼R	��w��i�P��ܯ�%=�����Jv8̳KZh�-�]L]�P�� u:v��7%c_M\B��J�j6�������y�P�O��䗥�%[LeݟrW��v�Zp�K.��
���Ǘ��6��~���;}Z�e�8~Z^��$����^��9ZIC�/�tu9�u���W~����ۧ��/��9��|�0"���AaD��k�	Ⱦ�:R����&�	Ⱦ�R�����*�	Ⱦ��F$ ��VS�����1'D�6/l�ⶣn�}�$�p��nG�,$��}��D�ߎ�YH��`�É�-����ۑ�-�{Zg!ٷ�'^��K�iq���8i�n:�-�{Zg!���q��qO��,����4N�8�iq�����f�iq<��8i��-�o'���B���YH��Ii�hq<��8i�&�-�Zg!��_�q���H��,��{4N�8iq���_�Ɖ�'�����H��,��;`4N�8iq���w�Ɖ�#-�����ю~hq���q��]'Z�hq���ǅƉw��;ޤ���YH��6h�hq���q��}'ZO�8�Bڿ'@�D����9�&kV;g�lM�1�<�ͺ���P!uE �{�AF$ ��dD�k�K&Ȉ����H@H]Ȉ����H@H]Ȉ����H@H]Ȉ��!��ya���j �-r�@('Z���PN��T��h��B9�"8P�r��p��D��@5ʉǁj 4���q���˿y	8-��@('Z��PN�8T��hq�B9��8P�r��q��D��@5ʉǁj Ԏ��8P�r��q����I�m���8P�r��q��D��@5ʉǁj �-��@('Z��PN�8T����8T��hq�B9��8P�r���6�iq�B9��8P�r��q��D��@5ʉǁj �-��@��-��@('Z��PN�8T��hq�B9�N7yǛ�8T��hq�B9��8P�r��q��D��@5z`N��@5ʉ�Y�@P]Q���rHf�.΋3CޒI�ۿ��u���"�+��2"!uE #�]�_2AF$ ��dDB�@F$ ��dDB�@F$ ��dDB�@F$ ������۴�T��h��B9�b7P�r�Eo��D��@5ʉ��j �-��@('Z��PN�8T��%-��@('^��K�iq�B9��8P�r��q��D��@5ʉǁj �-��@('Z��PN�8T�v�ǁj �-��@('�N
o+�ǁj �-��@('Z��PN�8T��hq�B9��8P�r��q��Ĥ�q��D��@5ʉǁj �oO��)N��@5ʉǁj �-��@('Z��PN�8T��hq�B�~hq�B9��8P�r��q��D��@5ʉw��;ޤ�q��D��@5ʉǁj �-��@('Z���sZ��PN�8Ϊ:�+�����O������w�^~�����������/�rP�
W���\]���\�
W��Ut�*�jpu*\�KP�5���թp-�KEר��W�µ�A*�v*�jpu*\K���kR�U��S�j_z]{]5�:��%��Ut���T�ڗAE�AEW�N��^�ct�
[��v�m��V�u)�.��t���q^*l�۽�\G[������k�u��q`*l�۽�_G[������a��Vǉ��u:l�w1t��qc*l����mu�
[��v7FG[W��������9X��e*l���]%mu|�
[��v�JG[�1�#1_�u|���e*l���8mu|�
[��v�OG[_������I��VǗ��u:l�w+u���e*l���Qmu|�
[��v�UG[_��������)L��e*l����cmu|�
[��v�ZG[_��������V�ZQ�\QǗ_t|�
[��v7_G[_�����{�h���T�:�{�mu|�
[��v������/Sa�t��+t���e*l�۽���QǗ��u:l�^":���2�N���EG[_�����{��h���T�:�{�m��$Sz�LǗE_u|�
[��v�����/Sa�t�t���e*l�۽����:�L���a�����VǗ��u:l��Z*�v:�L���a����VǗ��u:l�g:���2�N��ޫMG[_�����{��h���T�:�{�<m��|(����e��/�t|�
[��v�e����/Sa�t��=u���e*l�۽����:�L���a���T�6��2�N����SG[_�����{��h���Tغj��w�+�zT��ޫ��D]+�zT��\�{��
T>\��D]5�V�^���G%�����*�@�fG=*QW�սWA*7:�Q��jp��
*P��Q�J�U�ku�UP���zT��\�{��
Tnnԣu��Z�{T�rc������ޫh�c�j���9���Ra[�{��������]��L`���X/���W`����/���W`���X0���W`����0���W`���X1���W`����1���W`���X2���W`����2���W`�':�L�m}��X��:�L�m}��X��JGb:����i,S[_�¶��j,S[_�¶��j,S[_�¶��j,S[_�¶��j,S[_�¶��j,S[_�¶��j,S[_�¶��j,�2IǗ����� ��VǗ����� ��VǗ����� ��V�\QǗ�v3m�ej���T���^m�ej���T���^m�ej���T���^m�ej���T���^m�ej���T���^m�ej���T���^m�e�٠��T���^m�ej���T���^m�ej���T���^m�ej���T���^m�ej��*��/��f� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� �|3ZǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� ��V�͇�/��f� ��VǗ����� ��VǗ����� ��VǗ����� ��VǗ����� �쬤��T���^m�ej���T���^m�ej���jن�-.�dV_��83�-�4��v1��8�T�^�G�q��Z�JԵ��G%�����*�@��U�J�U�ku�UP���zT��\�{��
Tnvԣu��Z�{T�r�������ޫ�����D]5�V�^���G%�����*�@��F=*QW�սWA*76�Q��jp�f�:����)���X.���W`��*�.�U�ʹ�����Ra[�{������Ra[�{�����Sa[�{�����Sa[�{�����Sa[�{�����Sa[�{�����%Sa[�{�����-Sa[�{��y����T���^m�ej���T���^m�ej�t$���j��6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2���e*l�{�6�2+�t|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lm��u|Ym7�X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X�:�L�m}��X��:�L�m}��X��:�L�m}��X��:�L�m}��X��J������n��Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ��7�u|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lm��|����n��Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ�Lmu|�
��ޫ���J:�L�m}��X��:�L�m}��X��:�b;��Y����E���M��h&�ofN��lò-/���((��((���QP���d
���u��˙��3}g�:�v��8S�q��LbǙŞ3�=)sf�����/�o1�q��_L�o�!-��c�Bw�:A(�ʸ)MS?��s���n�fJ�5��v�e����r��G���Fc��+�@�&O�+j/{.J�0�s�Pn�L�ݺ$�5�+r���������2�3�A@(�\�����[_�hL��2�5uqs�_�{.�-�eZ:߹ٌa�;].f(���X���s�@(��%�u���s_ǹ\Q^V�)�)�w�/�=����I�d�d}�u�jV��-�c�,#�A��m7�}�L�v�N��<�<�>��_�mk7���Pn��ys}����v��v�%J���O۶f7���r˥���g_ \_����m��8m��/k��p�B��2�)�S�f�~��`�8�����E:��=���vq�Pn��b�-��I}\M��?vpf]���~��[�u�Pnu�Pnu�P�u���R�y1��x3�љn�cZ]I6D�^�^���ا�˂6��}��[*���wk�M�8}�>�DP�L�V�q
�\�}��X�Ɣ�Yg3���-�1!�[] �[] ����-�}�M�ZPr�M��?�BB�Ov��B��/��|AP�=I�_K�1�\f]�K�0m��>��8/�cB(��@(��@(���]W��0�%�E�q,Oc����'�`�a��� (��@(��e��~.9���>�����ǔ�g�C_�w� �~� (��A��eY�<�n5�K����i6S�]�љW`��P��r�����v�B�ݷ�Pn�� ��];�v�B�ݳ�fi�rf���3Ù��;�g��<c0�9|���pf���3C���Y|���ɭei3SJcY��do�q6��-y�'duBP�AP�APnu��]�9�������L�iZӲ�[��+����������2yt>f�Wrh�E��}���-Sq���.�r�K�����r
��&Wr�mZ̘�T���-.�e ��Pnu�Pnu�P�w������X��x���Ѓ�fs�f��+F�u@P�w��]إJc�Ι.��ijZ��X�=�0��<��� �T 
�K�ܻ�%n��)O���tv�}�sC�j���B�w�ʽ�FPnuْ��-kYY�c�ޝ++}Q�K�)��|�Pnu�Pnu�PnSD�>CL���m6KɡL��R���=��89;��&�r�!(�Y�r��#(��vkɹr.�j
J��Ba6�+y����[ ǄP�O��[u!��gB�5�ʭ�Pn�#�r�!�۹�p���Ù��; g���`0�|���p���Ù��; )sf��ȸ���n6[I���Vrv�`�ws(�Ű�y�r�P�{��������y��0��G9mf�5n͹������!���!�V�V��6�m/�,�|�c4c_�h7�mLy^�����j"(��@(��s6�)����4n&�����0ek�������r����;�q�F���5u�l����mYg��u����#(�NA��e
�wc.��<��қ<�ޤ-�ɏ}�P_ ����"(��@(�;��Cܫ��L,+��z7�<�ns���x� �{/���{Q�^�i��D�m�{E���1���9��mS���.�yP�uAP�=:�r�!�1�c��,��#�B�u�3aۆ���cF�r���A�_��[u!�[uÐ�n��r�⚼R	��w��i�P��ܯ�%=�����Jv8̳KZh�-�]L]�P�� u:v��7%c_M\B��J�j6�������y�P�O��䗥�%[LeݟrW��v�Zp�K.�����������?�������O��ӧ�o/��<�����//?-���_d��i���f�����JbW�ǩ�c�˜��˾`������@#���҆�,�c��uY���Ka�R������˟ک	���"�WL�O�L�O�&$�dl�j�{�/�Q��=~�JFm�
�}I�~� &e��@�����@p2��&��s�[)7�	�F�0�2w)���C��q,�4��ִl���;��=��+n���#���1�}\�pB+\�|���$_|�s��_�|=��M��	�^��&i����u�Ӱ�m^{ݼ�!6m>�8��%�+&����`Ю6��z�X�_���6g���C���{-F��/ʬ�!�}-]B�7�
x^�I}�l�:7=���x��W���G���2���?����Y;tӶ�.'i�x����p?�G��r����G����gY��hWt����Eo���;E��w�E���f�N�|SQ�K�8��ծf˖u�~q9K궱_�`ݎ0;�}pfu9�u�������2;�O�p�>��v�<�édΞgt8�6��X��?��lbP?S\���P�t�H5\�yB��+c &p����hE�8#�:�	ꓔN`���<~y]F�vLNP�t��}�>��vX��JifC�s��6$���I����#��;ҨT!�/:�9�wؚ��|aS_I������P�����!;Z��%�MwQ����8�.�E�� tu�u��Qtr_)��Q��H��,N��		$!a$p�[�"���ñ0;�c�q$/�"{q��9<;��f+�ط�5�f�^��	�'\�Cv�pN1P*���G.�^H'q�q�7+�O�D����:Fi�#�Y!S�D�	`�zc����fŎ�d��4��hO��d��5��Q�=wD���z��U�~�8��eoNj��I�x��mg8q
/u1N���ԏ�(Y�[:����X��{��������73�u3�-��es��	�a�����/�TC�.�N�1�˗�c���[���E��}ߙ����s�:¯�(������|#�.��I'�}^�n�Ii�?<�G3�i1~r�7����6���Ʌ9_��1�����|>��m��L�`�.L���_?�u�aٛ��[g�2&ϓ5>�m��n^���׿h�ҽ6#-��Ѳ�F�̸��흊��'�d��ンX��+2��}?�u�fΟ��nk?��!���O���7�4����;��	4Zz\q����ʄ�s�7�O��q�&$;OS�z?��|���H���p2�Fo��ݿ�:��nodf�滰�{����wh���TmD{'�x��½�}<��@�ѵ�W,�i�C~@X�����&�F�c@�:=���쏹I�8�����ԭ�_g3�%�(i�/@k4�O��C����n:��"�|��a������<�fL�dJr�v�nsȄ_?y3�u�jw�N8����Ϝ|�%w�I�-׾?f�\����g?��]�)��Xv;i�	�V�lx\��S�n���!�>���.W�lQ��������R�=�(�ˎb	��[���t�V��HC��*�O��4��*-�ٴ�\'J�<�Y�ه��A|�$��#�I�H�Px�#~$ԭLC��Q����"��T����3u�0tc��Y�M��59�P �6��ׯ��tg��>���η�s5wj鸇��Z:�x*��N0�x.�����T:A4w��T:��ϝ�Bu�US\��t0����D:��i4ЉL:�'(�Y� <�:w0�����Y�"<��Nf�s��0vv"����X�)R'�	�Ν�j�\��c���=N�`y,'LI./�aa:;�a�#��7n�e"#!�no�x�(���3��E7D�0�So��mtN�˵�>їЀ#X����=ԥ:��J���C�K-�Uܺr�bCG�C"�ô���;��� ��諕�a��AGh��r�Þ$#�nU��t�d�z��5+�mq9$��i/_��L��l��u�w���t�y�.�����־��N�5���.Z������弋i�Cr�C���㾻@���#��POt�p���y:^����y	� ��w�������>M�s� �,��-&��4�??� s�����u��&��%�8�f���n��ϋ�+#�8�����ZW��Y��@x^S���e Lu��0��(K8�3Q:�3�2�x��[���>�ĳ%���<��iT��H�6��/��K��]@�/Z$��٬?{ ep�z%�ಬ�[mƜ���=4�;��MI���@�29qL�xe ��.z��wQ��\�`�2ە�uep�л �@��ۂ�����iD��Os�ƭц�E��w��"������3�N��[���Ӈ���i��˧���}]^�_��_��?����Ӳ~�����/��d��+�v��&�sgb����q5}��8f��)�?W����_v6"F��>v�x%����_����|&���w�{r��w�	��_#>�T�_��p~x�2Nd�g�+�g�?����sݙ�C�E����,�'���	߽�9�hq؏JYϭ��%ݗ��c����qZ��R������I��]J�7ňX��OS���iM˖��Y�z��,���
L���%���k��T~�f�(�x�R��K�~���rO����rc�{�u��)�ώg�W�}|��=�u��)�o�.���x6�{�t��)�o�h\\i�Q�N�{u��)��(���W��g3.����!���V���P��[�:9�߹	똧a3ۼ�&�y3C�;3m>�8�ð�~߈��T��/z�����Mf���F�ۜ�g�}���R*9�<�u�iߊZB?�;��D����r��sI	)�SzV��_������ă���Ȕ��D�,��L_��<w�2��/������:ء���wo�4P���$\����)$����������T�dh��᪾���?J��z���M9p4])�I���^Nzkzʭa�`ܚ�w������<��u���\
������{� ��3,ie�{<��ir���K�ݡz�B#�k�{�����UBe	�6l�!�$�?y��;R����5�C+������H���'���\��vɏ�?�������W�K�YD�O���5�/M��N������-:\�ә@��G/�����^�,�6dB�w���ߒ�7Q�>ܸ�P��;o&�p������AF���̖�K eRS��{�/�55y������lk`�|��X�*0�
,�S����i���K:yj��?u����8):����*���
ciȌI{��I'��O}�I^g����*U�l���k�Ja�}\h5'�����u6܀�����"f+��7�Ux�#[��]�}��o�hE�p�Y3�b�������7gjS�w��}�dZ���^�z��2�F��p�!a�����tg�wpH���}��A����QX1�1�:F!�H?)D�B��y��=�-��~7F��L0�/vV��p�'�MW��"�x2��W���'��:s=�� 8���7���s��xpY��B.��=ݖ�+iK�P����3�I�x�g/l���ߕ�m�}�O8Qo;��<��m�}���г�x��lq�H8�>���?��Ł��m���Y��H��<+[�ω)���=�����_YpmN�EjШ�¢qUX�BVI�U���S�/�^.�z�V�;��(|m#�l`%���;b���+�������;,�Dg�g�ꝅ�V���x���I�(��J<�E��#�?������'s������i���{��f���]ql�s����m�Wv��Ǚ�G�K���2��M���Ly�Lr��q�����M���k�Ɠ��	��c@�����0��߲]Lt}o���LXF�ϹP\����H���ia���t2'�%��6��Vk��G3�i1~r�7?)��YI�s;߮���K���l���S��阒	c�Ѕi��G�lb�.�e(#�3q������6Lc7��pB�����8�2~[SY��&tf\���mt9ei}dd̟EL�"8���Yɨ��J�)�����8�Ɖ�U�[���a0CH��cJf����ӜC׏[��IĬ�$ܑ�]�T�.;w��i49nބd�i�S�Gq����o�E��D8����y����&��+9V�����:�.E���	DZ0C������n�n���5: ɶ���*����:ݢ��[�Y�����9�cMc�V�
+��
�4������Nݚ�u6S_R��u��FS���:�����z���j��g��+�@V3�e2%ɝ���m�G��a	�Bz�A;�v�H�m�$[l��M�mQ"��w�\I3��g?���\Z���m�7�5a�J^�m��5{�m[^��_E">��$h��l�
�'H�B�;A����t��B��� �7H$��R/J!q�@/�!NV/�˒HH�(���/�;��˒�Τ{V�]�]�o��)=j� ݐ�3VQ��������JbC��!�!����(E	�預��/
	��߰/@!!�䌧CX�#����N7���L��s�|8�۱_�G%""}��5S�UO>�x���|�m ����\��o�������'jT�yX�QX Y�R"��Xi�2�"VZCΪD��*Sd��#��X�l:�h����*���ڏw�I�G`Y���. ̛Y�q�D�w��^&���9Ъ-�/��f�t��Z�]�A�{g_�#�};��G���^���>ݩp��+����m^���]v9'��:)}K^�����<��*�V�������:���d�j�l����9�F�6���-{ǵ��Ux|U�(��	Y.���J��-�?������7���p��)��W��cy�xVg}�����(��5Xų����	�r@��ٶ��H��'����XE&��W!Q���x�ƼY`0V�:k��W�*3��=FD���F<^C��~�V�v���;�W�,��������\1X�++~r��*�Y�:�:ϟ�#�G�
VQ�� �gY��_�[@r��xO�;���go�kO���#�6.6��j�wW�������w�[^sa@=�c+��yB(� �R�GW�	a�!Zw�]�'���v�̷��}gTߋ��y�;K�w���2��O���'T�#�c	r���o����`O.<7tnK�o57�v�e;\�U�?���V��{���=XB�Q2eőF���v<Ja%<�9}MX�J�@?�sX9���s����������l���%G�{	��Z6��T�5$YЫ�x�LbŬA����E�y��(.dU���P�Ad%ܞ��<�w(��r����ߡ���J����m��������q�
y[\ɬ~���.�yK&�n�]��:�{�9k������8��E������
��cG��}	���íW����o�-Y|�5�B�"�WE=��<k�����f���X�u��ؗ�����c�����NI���7���z����It|`9O�x�ۂ��8i�RDL�Q$�?*�S�h��o͟�D��<�G{p��g�0>�ءz/E��3kݺ�S��&���Eq��8L����o��o�?�d,�p'�����(��~|(�����,_D�����Ql$c��~<�S�_C�Le�yH�\7���3��H'T�]��"$E�\(qD<G��H��;�#ħ&�Y�ڽ����Id}'�/s�QO�P�x����#k�ȟ���O!"�(���/�0��gz�WE� _��V���:�L�W�?F�-�Pq�����2��Z#&r���D8�ם4��r�%.>с�lK��E%rY�[#U���ȏH;V'���%�j�x�}k��DN#+Z�y�<�(� kͷ��j�(�5�T�)b��~��KS��6���eؿ���Ǘ��6��~��������#/�}|������ßD?�T��W��4�B?�T_$E�gR��S>!Z�g����<!J?�+.H!�+��u�>�����n
�zF<]�A��3G�g̞�Ѿ�g��O�=q}�Ծ����~F����9
?'��(�(�}�O3e���O��{���Ws O��Q�ϡ_���� Z4_�Cő[��Z6����T�(��ձӔWH)��eC��tZ+�t�'��0ǟ�q{�ާF(˃%F���� �������N��м��ey��� R���g!͌ �χ^�pI8����R�|�1^Ϟn����2B�����0^O��&��w@ʾH�Z%K���AzO�3|�?<��B��`��̝m��#l��1^+a�n�0�=�Y��W4�j\Bxv	Q�@��,V�==�l����CH�Ӄ�&��ad>��n8�Lx>�v?�|�yB�z)��Q|��v/�y�[��� ���ey΅�� R�	�~�V��t.�R- ��G�9�k����CD¶R<���D�r��2f9��QG�r��3v9Bj�v��v�\��!y�8r���v�y�kG�r�ׯ��y�1
B<�c�x*ǰ/�O��!��1
B<�� k��$���oTBb{Yф�D���Z��ZV9���	�����Z�к`9��e	m3$gq�(�,�o�HBb��z#!1��"i�bD��}�Nؼ� 2Kk�	��=��t2%Db�����HL� R���e��a#�Z�}P��E/�ܔ�_��||�D���!)����N�^�����A�O>���
|��A
��yFNMH�=!��c����<��A�Nu�\�#������N�jv���#D��"�xϐ�W�<!w�c|���lB���Ay6?!R���>�� =�#Hᛐ�����:b��9�j�d)K�K d��8Y�a�E��G��9=��q<>��VJ���ozi�%B�?(���(	�㰤Fj� ��
� y:�H�~_<��Q�����N�/KzPZ�(/Ǹ��Ay�����%{1�,��[ް��� $��\렴a�;x�W?��l�F� R��\V場�ú4��,�Ai��e�ʃ�/�tP��}Y��� ��"�����rY��� �ȋtn
}��W�����ׅ>h3@9��ׅ>h�h91�u���P��j�C�o�Y\-K 1�u��Bq]��C\��,������.#�2���:?(�I���C�0�j�e'�!�^�ݠ<A��v�F�4�D-�ojwPZ�8|Yh��O~z�϶5QZ��,ǰץ4xW�'yD��?W�Hi12]F�K���3(B𽬝Ay��e��'�i�
?4t�$�EH�/�aP���	�W�qS4�� D�˂��O�V���Р�����%	?oqTR#�l.{נ����YM~!岆�E�r{]҂� ��˲��*O�Xt�o�bPZ��|Y�� ���:t#��)qY��� ���J�!�,KAy0�y�[�]�v�����ú�4�?�ö���&�ǐ؛��\��@J���\|(�� ��hE�{z )]}jX�;�Ge1��rYÂ�"��u0(�p�p��8�c�R��:�!ž�CAy�;.�PP�����Aȩ/�P�aBN}Y��� ���:��Z�_?�}�d>�?���׏?��~��?��Q�~Y�U������-�\�Y?.?����4��o��_�'��o�F�\���Y�@��O�nO��S�d9#YN.?G�W��~Y?.?G�W��~����#�/=Y�����#�/��_&��������@�o ��������Qv�Ͷ+d���p�tekH�,t��e���5�&���б�5�l���3��v��
���c2C�f��r�5d��g�[��ϑ��|M؉��Q��c���z�,e[2C�f���֐mg�����[C��!3t��f^�g�����r�� �L��*��<�my�����[C��!3tl���;7��ȡ|�ϑ�my�����Ӓmy����[C��!3tl���^l٦���0|H��P���O�!��;6aw@X� ��x��!3tl����lٖ��б��>�$BB��:τ��I�'�=��;`�� ����
*[R��!3tl���l�%hl�����i�P��	O��!�j:��; ,U����:6��k��lDf�����o�"Q����Iٖ��p��=-ٖ���0|X��筁���:6ý� Y�ȶ<d���ô�B�(�������3a�l���б�M+����c3�n��E��A��&��D��l����ᦋ|�c���%e; 2C�f�weakȶ<d���po!�֐my�������!��:6ý�YÎ�q������!�X��б��]��c3��.�5d�2C�f���bkȶ-d���pow�֐�C��D��S:�O��>��б�m���}
��c3�[��5d�2C�f��wck��)d���poMG�0�}
��c3���5d�2C�f�������9��v���Q=�_E��z<�~�#T�Gя��١�za�_�Gя˯��!x��ůǣ���Wѿ�^����Q����_�~����я������_X�Gя˯�!x����ǣ���Wѿ�^����Q����_^/l���(�q�U�/D�]����/ۂ���/l �hH�!l�wl �hȶ"��ު��^9E`{�; � ۝���/l �h�v(���ٻw�l������YT�����
�]��d��!3��_� x8-��G`[��!� �����Kf�2Úv���箝aw��)�EͶ<xw@t��my�k�6 r4d[�g����hU�~C?��ưOc���ٖ�̰�a�у��ޚB`; ��!� �����Kf{2Úv���箝aw��)� ����Q��̰�a GC��yf�0-Ϛy�
�-�,U�my���9�)l�CfXӿ���!���4,l �h�65d�5 9ҫ�nv"�PӰ��#)�Ԑ�t(l �h�65����N:-�o�*��8d�G�����G;� ���Q�oX�^2���t(l �h�65d�5
 9��lSsסЊ�OM��@��l�CfXӒ���!��<3|���چ���Iٖ���C!��!�����[6 r4d{2Ú��٦�̰�a GC��!3��A� �ѐ�b�kz6 r4d�2Ú���w6�.�̰�a GC�m!3<�A����q��lCfXӒ���!۶<3|�E���_�!aa5�pM�BTz� z� z� ����6 r4d�2Ú���٦�̰�aa GC��!3�iX� �ѐmj�k6 r��M�aM��@��lSCfx԰��ѐ�bp�!o��!���8/�yK&�n�]��:�/-	���*Z��Q��z<�~\~-	���z<�~\~-	��-~=E?.�����������_EKB�za�^�Gя˯�%!x��q�ǣ���Wђ�^ش��Q���hI^/l���(�q�U�$�6��x���*Z��.ۀ��Ќ�mA�kZ6 r4�����5 r4d[2Ú���v�̰�a GC�%!3�i:� �ѐmK�k�6 r4d[2Ú.�����̰��` GC�E!3�i+� �ѐmS�k�6 rv��>�̰��` GC�O!3�i� �ѐ~d��)x[�@��l�BfX�8���!ۧ��t
l �h��)d�5� 9�}
�aMk�@��l�BfX����!ۧ���l �h��)d�5�  9!l�BfX����!ۧ���l �h��)d�5�  9�˻�>o�� �ѐ�S�k��5 r4d�2Ún���k[�$7����Co�}�,)B�6$����`�ZZ���xm+�A���.��p���)y�3;de��S��DX�`��SKx�i+l���qJc	�9�oE�mt�:Ni,�9���h��[�)�%<�x����n�4����V4�F�����s�ߊ��u��X�s�[�`��SKx�~+l���[QZ�)���V4�F�����s�ߊ��u��X�s�[�`��SKx�~+l���qJc	�9�oE�mt�:Ni,�9��h����qJc	�9�oE�mt�:Ni,a� ����a�8����ط��6:l�4��#�V4�F�����s&ߊ������q
�Ļ��a�8����ɷ��6:l�4��3�V4�F�����s&ߊ��u��X�s��[�`��DZ�)�%<�L���a�8����ɷ��6:l���p������t�t<|�$�yN����dО��R1��V�J~^�/*�e%���ו����V�Z�T�����������������������"��(�(���t�wD2>�FN�G�x'�P�� �_� �uߛ�#�Q���$I�;J�Ohw�єޏ�/��Kʧ�JBݤ`v�؞*��fWsn_z?�����3��Q6N�g��N��	�&!�a��1���~c���y�w�#�<u�Vr�,<J�G��?����c�Dw entO$�J�ޏ�/���So�U��4��v������a�8������Lѵ��)���L�/�N�cW|?���~KUo���L
Əy�/�ωk�.��������/�_��)�����A���O�ڕޏ�/�_�a�Vf@N���^����h��F�ޏ�/��m��Z�;�o�vN���%Ƶ-��_�����/�?�L^N�FND�����irv��(�J�G����/��_꿷��&�H$���A2�&#��`R���c�K������/y�NuFkSG��~r�_^�d�$:K����(���a�K�����n J�xߏ�?ԑ�B����٢���/��_�?��4�b�����Vb)��[ezڹ����/�?��4����m��L�=���ֈ�}G�7���0�����/��_�?����xN�#�@]ߏ4Q=x���������/���B�Q���w�`�:�!~����@�q�3`>M��E���_�����б�t��Q`:�~ �0�0p燩8���K����m�� !��/��P��,���B�r@8�T���l$��Z����jQX�F���a)�k���l$��j[X��R6r4�M0��^�fS���TF���h��˳���I�B�A�aM�����)5=�q2^��a�������G���������7ɕ$v(r!�FD�h�_ʆ`�K���ZN�j��3�|?�N�B�^/G�l�D����/��_���;�z���M��M:*�g�Zn׺c�K�0��c����	�Q���#��~�z
Q��e���D��!�b6�_�G���o��lB�$���S�Ntt�����K� ��b����sGaրyT��T�N�u��L	-������G����/8Q(�����?��"ނ�!2���I�����/�����/�OM�X��v�/�	��
foχ�Ӣ���/��`��C��?!B�� !B�� (�Z���q\��E���?�jګ�d)8�5P�Rp�k�����@-0K�9��j�XkK�9D��j ��R ̳�9�9��nt�T=���c�K�9���i�D�^7�z�=�%l�"�m�9E�J%0������g����P�~���$�7���s*������K�b�B�Q�����:ϥ$ۀK�;O,7���R:(V\���j0���)8�:�1M�'�3�zk	��4P>L�*�(�Rp��/��B�{�9�,h�N����@p?p���=�Ҭ�T��/�
b��G񗒳�['�R��Az�zb��y6�j�E���K���\a�K��3#�O?�Pj�=��~?h���E_,UA�K%���c�K�%���C�N�P#G��L��1���ΖK�0����_�?1�����N��w�0� '͉�`�g����i_,UE��p{����'7�ǉh
��J˾X���/�*P�|g���� O<7�����W,�D�����/�f��*�N�r!�iX�T�����}�z�o��o��ǫo�z������OW�1)�?�H�����?�X��͎0P�@�-�,P�@�=,p���wm��W ������#L���4��S�~Ā)>?��Z��Q�}Ā��>b�P1`*��0%�1b�S[�fD�&1՜IFLd�����$#��.Ɉ�XK�Q�dĔ����,�'��Y�N2b�����u�4.��/��J^^�%�$#f�g����0����,3&3���䫒��$z���I�4 Ri�!b�$#&�M#D�fD�?Y�a|�,3�q?�q1��1�5>������_��ػ�)x�7�0���O��s��n�ﻇ�f�vf
��
�hY�7�ݣ���Inں:p��P����˧��ɍ
����|�R>Q'��ظX>S9��J��B���J�+%�'t�D���P��	�x��*eR	���V�()B�}�ẝ:�lB�j��+����І+�d�	�l��u2�@�*e�N&���Lh�����P�PU2�K�2�Z�ZEɔP�Ӌ��"s^m�*a�v��ڨZ{�S8�� 9�tQ�	�ךQn�$\�[I(�X��I(k-��u^���X�Z3"�B���X�Z�"�p_#KXk`D�(/o��%�vg��M|�t,am�+#N~*&�u��V�C�AKX�d��9%�S�F��0S��Յ@��%f�:���IV�$冋:�.���&������K�:�W9z������ksr�'��fh�����"���R���u�x�����*�b�ԋ��DU.��R/�:�R��Tڌ�Jt-������ŎE]R�U�1�=����R�Le�1��2͆��p�=%,�|��Z)��iOٴ;
�F�\4��E��(���橑0��'�0�cߐ[wD�Z8�9"G	7m�KH�u���&2���ˉ��
u��Z��oy����})�I�|	��Ԙ���<��C�0�aߐK���OI��Ґo`�NId�ٰo��S�)	��UsJ�?%a��G�Z,�`��W��L5�1ҋ�*v �ʆRX�*[v��Nc(a՞[�D���Bx���Z�n>~��uL��ӱ�}�矤����,�.��}Iw�P4���Y�}�u�P	�Xggzd��")��	���;V�*L���B����~$�La�v
���
�H���Y3[��*ej'*�˧c�J$�Mm���4����:;�[����)L��9*[���H=!T�4SX��
��S�΢*�×X�1u����
��{L֢c�^�%��I�Zt���j*a<M�E/Ttb�\b�3u�`�B%L����U�Τ�B�&�;�$,����G+:�w%=M��t��O�-������~3=�$�q�H�����?��#�d�G���£�����L��������ױ��f)Y,&���⎳��,�����3?s�3=�s�y����j�g4~6���}��x�3>�����s�x�?>��:�s�y�w1�O���sd�9�A�}�/،� �>ȸr� g��/r�'籕�����q�b�'����b�'�����r�XN1�L�8��x���?��߬3���,��e�/z�U=�)c1�3Ì�|*�ɸE�b��Gs��ѹkq���.�L��T��,��%Qs�T�75kRŪT3�T�0�b�c��a*F��Ѡb4�Yc*V��U�b��Y/:֋���c���:u�c��Y/:֋���c��y/֋���c��Y/:֋���c��Y/&֋��g���Yg&֙�ufb��Y/&֋��bb��Y/&֋yqb��Y/&֋��bb��Y/6֋��n��Yg����O�n���;����)xo��&!�����X�%q\k�h�)D�V���/��^����3�T��s),�P1 oM�4ieF��^ᮥ;���F��V��O�
�u8��iu:�W/� ����-w�u��ܶc��P*����w��Q�:�m[k���ж������߇�P��ks���s&̢սt� �9����ZCיJv=����׬���ǟwO�L���~��������v�����T��S�),����_�Ox��~> �p�ݧ/�й��~��M_���������w�/���	$�p�0���ۇi����w�ݟá%���9����Ͱ�������d��{��U"�S������}8��OW���~E����v?����_�?ҟe��O��� �o���O?����Ϻ��(ߒ�UJy$���>h��A���������Zf��X�,�ׂI����04���pe�WҤ�:A��Q�S�!/�젺���qzxܽ�}���{�]C��Ԡ���J�,����s�0|��p}0�*.�1��������g�}�k�/�O��2�޿zŮŵ������`n�"��k�9�P�)A��ܨS����%�p��^����� �Ƒ��nq͔5L+p��ۨ���Nv��G��żjd����Yws����:ekßw��lg�����g�����v{nUʜ�km�����F�8�[Γ�Ǹ���]۾4������.��B9�#�Μ�u��N9�1k��g�/�:x��]�hi,�>��.���_�!�N�k�^�K�e.�u�i��[��2�A��%t�tIg0�}�
�����#HX�[�&S�w�T��c�� E�����7�'#[j�0T2��!�&���D���"NO��p��^�)��Q� fh'NcbF]Z�,�����`���Y���bC������S�h2��$tXB�y�&����W�m2H��0�}G��D�@�3J��_Q�,��b�M���uaHJ��($I!I�8�bpRn1:!#�ŧ���e�}K���-M[�4]l�b��2괓�����1@F��-rNW�1�2�\���\ƶ��oZ78)k��$��O�f��m{/�AW����c�Av�;���)�:\t����!'�z�!ٕ��>������ݟ_�0<}�����iy����}y��x�x��,�~���nx��0=�D8${����������]Q΍��Z�<͔|�a���>���
�N���F
��UDy	F�������P�e"�)E�Q�~�����~�����֗?�*rt{��,�w�B�	���=�����;�J���i?����}�c�,����|��9�}��Q�N<��u��	:F��~��T��¸'�X5�X�i���ec4dcxec�f� CQ�TB$"|�h�!<�V�`<�0}m%�VH�v��n8���z�����1ݢ��ݥ��> ��a��;��ke8S�~ig�6+F����3,��?A�^��5�?�튍���RS%��
܂M���|Y.��Db7G����_��4���mrӨ��1�5����V-����r�\���4��0h�0�|�0x���@��='��7I���G�l�E��f�0�(jyo�ts�e��}\u����d2=!�>�CD���CIv�sl*�݃�8M7Gϯav�n��q{��9��'��}�c���eޛ���������K�9M�[�.�A�.�U�.�i�.�}�.���t��2�k�����>ޖ��<9�e��������q
�g���G-���je�R��:x摣�G�flPk��{ť�q�8b"�O�m ������x��=�T�	����XF��)Y�D'2�-�=�6���e�D-'a���#�Ck��=�����Q3�*`؃?�����z���fl�K��s��::��H݇s5 ��̂�f��^	��>c���"��s���(�q�;u��1���#`T��q2�ZR1p�x�')Y��}vE5�g���\��bÒ�J���h܌�3�;�(U��c��$sJ҉�������eD�����H:G�i:�xo���3��������юRN�wB�D;��P������.=���k���4�b����B���Pn���j^ЇO�����8���0�M�6�~��d�`�HCG0��e���Sb�J�d��u_z�z�7'�g|3�<�Ŏx���e���@<X�:8�!�"���/�F���enQص�y���K�/O���>a����:w)�J�':�!lN��C�3Q�&k����㌳5=Ao�Z��'4�Z�2\��]>ʹ�FC5���!���$����S��0������u@{�����O�r��z+]��:ϥ$���3�;O,8b���R:�Ω\�U?�&�Uﵖ���'�W�F���z+�Ү�Ӕ�q���񜵄�q(�^����W��m⫞�����n�[�.��^x�:h�XL5��N����Q��6�0crz26�u�}B7�-�p;mB�e�[�����{Nz�zb��y6�j�(+��;����O.�~⼡���_��V^��{gF���hC!����Q���V�=��yRٻ/�Ie��=G��˳�j��';9tB�d5��2��aDx� ���8�Ѩ�����'�����:?���_]��r��WFe�ЗG��Gv���(�:7��(��_�U;s&g���_���d���E����^�������o�����d�Eك&ټ���;�敹���6-_��M鉓��.�,MJ��8�?Mq��4A��4݁��Ó&8�$���I<�-~�^
���1�k�D���IS˜���:=*�9��@r��jjhg����i
�̾=gіR��?{��r�� ��0��
"H62O���Hj��Zi��¤]�!o,2�G�W�j2�u(Z�!��ND�B�A<����:�p������Ӗ^�P;��8���BJ�[%��ʅ�����Mm�P[��N�����<���+�/����6@����v|��*�H6�a�/��v��7WZ�R����Ð���4���j�o������������`�׏��O����x�O̺���x��������ۻ_��G��Qw���ko����m����]�ݏ�?)-y���=�=tn�ۉ����������]�����U�y���������c��7
��J_W�w��iB&Ԃ�}�� gs����E �#�B )����hda�J#`Ag5 ����y[ �� �Z�Yg; �� H�~6  :k���b�ް��]h�5�R�݉ߘ� "�N��n}K�{Q{$�?�#�10���Y��^��0�� ��n���wɎ{���' �t��v'��	Ӄ��o��t���~�c�hZ��Z�/��G�:c�I�4:(U^���hk��t;|�_��6l����(T|!4*���pU����6E��ۡ�n"�ׂ�`A�����$8�w�L��!������!��kg ��=E���F�,�Ĕl��B��pۡ�d0R�����0=��<�9���}c�� b7�n"�Ud�ޛڳAėc��lbB�qr�mH�8��3E���1�LS�C%���Z�"�(�	3�X�-	�(���kq�����v8n-�Ga��5tX��7F�k��f�!��ZE�ICa� �5txKd�cH�DG�Hl�� ���ol7� 2Q<������l=��R�Ǌ�6�b�nЅZ7��t�q���=�nl]��2 ��6��fP�{��N�i�G�E	8�k+F�:�emӮ�m7��n8�l��Qj�K���r�7)��5��Q�B�]|.JlYٕ�����Tf]��|x��lO�֕�m�R���q��R�2�A��\7b���a�R��to�Ѳ������]�����
��L���ް B������[R^��L�\	l#��H1ȵ��[v�I�lY���P�<Y��F�sA�,I��޴U��/Bs��� H	�!q ������Ӂ��b�� %�� �
M3 Xҽ�%h���.e	N����HY��a-�& �m7����Mڽ�����hT����tBh�u�]j��^AJ�ʬC�,��p�*m���]
L)�k�y[�$���t���Y%ָ�j��� ��W+W���k:Mgp�1��m�˖c�N�J������t��|n�Ih`�Td��E�:-K����v�'�Ǌ�g���t�r_�MbH/4"�y���v�Q���w�	��Xҥ�A!$�j�����W��ن�qA�!��Y�h?cBK���ղ�K��B��L��jY}�6��I7�]�Z $��t���=X:4������8�.f;���K��$!\1�r�K��6e;� jE5å�z��ز�~mu��1��pdo[��r����QPA��R�rM-�C
�;BJ�zh�2�� w{������ȹ��*�%)f���:{�r�>�p�	H����V�/�-��q5��)X2��ҏ�p�1����t; �D��������$��#2$�&��o�ۍ5=[�m��	$�0�k$�hI�A.T�Ȑ B����y\|���I�]�V�:?��τ��Ď�M>�谧�nrlrӪuhN]��d)O-K���j=�0m����M�Ҵ���c*/�.�#%%|m[��ay�&�n�ø�T'zJ&:X"�@�ER���Ӟ�ɰ1��H�������/��^!|�٬F"��[$WP�7
9����v/�[�
�kOeV.�%�&%�؎#/gA7W;m�_��x���~����,���t �e���.4ȓ�m�?��q���MK�7�^�F�����&��ڃ��MM��@��{S�R�|=
u!��I�6m	�1��xS����g�/j�����'�%ݛ���j���#�>Y��� H	6(n:��WyS �WA7w)�\dm#��5=��%��B Y��n�R8���
�υ E�Q�[B�!+���]��F�6[�ePX��-Z�
Cs���ɵ�6��PATa��h�`����)�υ��A`���+M� =Z��tŀ�S�[!|��u ����R�;a��6�8� ]�U;藅����%�b�K9r'�y�f�O�gW�i�N����W�DFLv�!/&
W4���-�vC.�^�L�e�<���#+��ͭ�a?0��v������3e�#��Ըc�Y�6W}:~��{~)�k���~�i!�ߓ�<J�ܪ��hQ��k/�X&~2b�"|[�e���S�.����B�J�B>�uX���qh���]��o0����\R�@`�S
I����ͭ�Q��v��ʛ�������g�<2Y5��Mt���Y��ġ�rq�k�6P%e7ué�.����僚�5yӃ��ծ'R:C:����xχ��iNX�7�h9O�:a�cΗYd�d��:���,�t�^��&GwA�0��8����������+J������I�c��k���f�m�(�mAt�B��kf��7b��m�k�آ�U�O��b�Ft�����"�pБ7�b���l��[Y� ��A��v��f��2P��!����ӑZ��ˈlN�Ic�E��"(�rZ1
eb�#�� ˠK�>�)�b�#��¨5犠E���(�D8ӥ��r�I��c#з�b3J��=�ͭrpѢ� Z�u��,o5���yH2�>F":nM��q�ث�9䜇�Wt��9-�J�-�P�����H2����3��tH���r=�FZ�ed��22_s�Z�uH[�s��8�K�GN����C[�n�{��Dn��5��E�Ъ�<�xyGS�\1���)��Wn%k��ډ#KW�Բ��9��⤖�5Q|�A&��fr��6�K���(�g������t��f���(o�%&��^�ٴO��r'-�������DM��l�|�0�V盢ddD1�M/O,�Hh:$���@�
�#�tu���Y�iw��v Z�o�L�,QLg2�E�M��DFv賐����f�ia�e�.6C˽r:s'��i:��h˕t�Um�ɶ�D-�O؆��c���];����t�+V��W4D�{�>��"3���X��E�Dfmi��ĉ\i��ȉt����"$D�QF�Cr����I5�E�Dz�t�<�&7��<�fu��֞���D�6�눖��|��6�`��r�A�u�"���F�A�<5���d]�AG��X�m��e�o7�kK@��3�=�K:�L�%��t��
��e���;2-WV��hQ�Z�Z�G{۲g(.�Tz�`y��	"O�g]c5�]�2Ìu;��0/w��N[Y��}Y�������|2Ö�c�bCfU�<Z�u�˸8slג,c]�e?h����p��~��[���iz��>=^}P����������ݗ���������c��wy���m�~>=���n����o�PK   ��X1	���  t  /   images/4a240ba9-1e57-4d57-96d9-193d1ad0babb.png�x�_S۳vQE�.UzQ!t���J��C�"P�# R��"]�N(B('�"B�H�;����~������ڳf�<3k�<�����勷/�@�˪*�� �Ym�y��y��]��猇��<���q���iȁ@屗��Ɣ�*� �'��̤b�TU�Ӈ��M�f�d4����od&�]���E���N�����/_C�������O�+J������W���/�_��Q���!7����ʺ���a߲G����K�z�b�쁪�/L�z��O�yֺd�ݽ�"����J��}��~�3 Ѓ'%jy#5#�թ�GkF%�x/��K�*��y�R��S3�VD��r���v�!�>�'�`���沆=2M�5_o�A��"�����b��3M��iXMJG�x��i����P���t�p{16��C@@�m��
����%j��@�A��!ax�贴��<����
.P�����8TC*��yk?�+����ز�_��1i�)����~����ḣ}�t�����C�g��������{��jj��ks#$�?�-,��TpV�R X7���.�\C�iX��C�%���S����V�S��s*�z��ՠ[�q��8�mM������cFlx�&�9�07�흚�i^�XުR��\��쐰!�\ܜV�ϼ1_ΐ\�/p�y/�e��jv6��i���E47��>���"**�w���2�#^��q�ˆ\��7�e����E�Gz�<�9���|[f,��	U凝j�fceJi�e�>^�c�G�s(&��\�L����bn�jﴂ��5��$��;o)AGq����:D|��yg��N��<F�����+T�bP: u�볌O!���[���@6�V̮������?{0�ͤ�?�q�E�::B��؏���K/��ED��9"o�t��i��a�w+�+n���Nc�!�R��]-�Wk�O�KW���P�Q����$��"$/a��B�p�E:�������,�9�EL;���8��3��R��>8�o-PT������g-��>�4ufo�]��:�*�����GRd�\�ʛ�-HUߗ0
P(g���"Q�ڜ��x�2���\i�8�Z�g.�-���m) y�2.��Qov�~�*	��nʯ��t�����`�g�~C�'
@��x�>4O}�>����:�pU)�#��t�Z�q˹�u�m�l��\�hK2C���$%-��W�&R�j>T�JM@��m��!cX疩!AZ�J�/9z�ޙ5o��nn�Ñ�!�.���g�
�.t� P$�nx[T��F���2�EJ(ڭ%z&ۼUj#Y��H �0w���{|�b�bzv�GX?��b3��+�E�A���E�e:r��ID���Eok7�3��D�B I�0ns����x�?p%F�HiC64	�Yƥn޴Ο0��b���L땄0��-�	4E�Dr���#��۪�k�ISp6�_�=��+;�0��o���'��Q�i�LA�!�n�/������/.E�V������٠g�@H��\��2�Q����T��Y,?���j�:h�fh���&d>���ւ���{_<%��aWx@9���8�����ֽ6b���E0h�Ѻ����Ubи�e?�8��{�S,^�[�32�p_�,��4/j��Y_�����؏��W����e�ax��}����a��@���������V�8��/&`�I�~5�X���($g ��s��٤cʧ�.Q�Vw��LÜm25�w��i�!� j���(k)�,C�ט	[�.h[m��"_�F>z���Z����/?`�m�?9�-X^���d�Ve`���:����)�}��`K���w��m5?l����~�ɖ��b���
v��'"& ��" ��O�}��5����B?����PH�ି�FQ�#�[�yh
�!�'�q�1�ޢ���T����	e��\u��&��0(��.�'3�b��q�H�c��ɲE��}����2
�7~��f _L����	u]�3]��ZI��Z:z��ơ����m����{dpm�OK.π�	�U�`0yn����!FG3s=�v#<0X�n�p���Cn��EVKu����7�걾�U�y�5z���^�������������>i�|f\��.C%_����v;j�YW��� �CF	�����]&������)�X�x��5���Ţ�oA��ɶ��������qXq����r��'��Mk9�K�{�%(�~��u��B�y�b�q�4��;!��;`�1ʎ�%q��:tˎ=Y6lF�p�[�]���j��/�ټt1=�r\�q��=��@��N��k7w�E�֊���  �~��*E�/����)�>,�!~)d�s�u诞�x��v�����$*���[�����W�j�ɀ��FQ�/#:π��o�G*J�^c�g9�9���D���Jy�|�z��P�	x�^Y��j�� 
�B�m�Z��n���R@�� ��w��3��� �y�^�N���
�ǋ����%�( �H�:���On����!L@ ���\���ٷ���ܮO���k��>��\���Z���N�(短��,|�,�%`�"5	��~q����{!�m���e��=���D�na���/�
?���U��ڐ?k���U$a��5	�f��EI��7~[)�@W}��_��Z��z�����{�짨P�*���J�j#p�h޷+!�7������*�qK�ʮ��]�]��M�.�_W{ˈ�m���N&VW�JMM�~6�O甤~]",�T1ͯ�K�xj���߫6?��߫q�嬜��J�G�H������o���t��я���I�N�J��Ŕ"r�ҥ�B��0�90�la��#3��C߉��2�����e�޽���U�58��$45W��T�i"��5����{���wYY����"��W6�OOo���S����UU�\\\=��ҥ\�O���[':X���WW0�����X��b�<�?w(��d`
�%4�&���j]��{�=�:�{(-^�>��zz*xgc����!���h�sI[A��@|���N���/s TY�̙mFD\\��}� ��t�� �Z�/D�,��#���(���i)��va�/�/t,�3$&Fio=��9�j7����a�e,�ګ������^�=�Z�e
�A?���@��>H+;�X̖��o���rX�1����p�0�ڨ�V��8hDo����uޘ��9�|�2���GNӞh�yV�lD!g���)7��)����0�޾ޢ:CpOo!��P��.�~���6T+���v��ju�:y������L�"�#��T��^qf�7m��<�-4;,:�/1ʔ.,."/�^wpO��7�
�Ʒ�w���H�P�Ÿ�R<�\[J�Ú<�@,��e5si�4q����/�\��|�؄ؘ$0�.Ӽ�Se����Y�S۴F��v7�e�3���h��|k�ӹZ��ַ�a����_&��=������2��F���}u��k�O���ģң�m$z�#���.Q��Ӊ��f �>�'�$d��槻?�P,\9�k�W��3 KW�s��V��y&���^Ɍ���K��Ɠ5�G֑�����K�(x��vu*u����'�nq_�W�3���&|Y/L��b>��!�jM0���6�3�9�8m�q��v�YY�6�b0�i�]��<���IB/í�.��M⹬��B|n���6<7��6K���e�A�Czt��|�V���H�Z�U}E�]��D����]q�
=����Q%y��J�]����;�(�fEY�%�W��}��G�߆�v]i2�Ҕ\�ԛJW��s�R����՘�4�ϥ�c��=DS���>��N�Ni�HN�[��pU"m�sP�|�8	���8v�b��G�]������	K�W.+�|5<D'�^�0��&�Q���@-
�P�~ �^޶Fi�(6QW:Q��ca��	F�C8�\S���ہԲ2Ox�5f(�L]�A�_E2��1���(��do-c�X�Q#���"��F�V���vK�n.�Vv)��Z���f�>�Qc�Tl�-��R���_}��lk�7���W��MY�a���|`'yH��y.��y�+�>��֍�$%3��l�[�$+ݼ�H��)�+e</N�-�]�j�fn��d7e��w ��T�
}���׏zLG�d����-�}��N�K�~!�r#f�\��|-�0�����I���K����Y@�W0q���iPzg'3��0d��HMs;
�J���^ρ�pn���C����Ԏ�̴`�]Yk^�j�������N��/��O��?�c�iĔ-�o�rʙ���U�HVT߉<�O����}.���I[�U$�/�0�u��d.�,,"򼴈�H{A>���l�K�u�Y`^H3�B�,>�uǷ ��Y5)�dB���X8 Х��er�ԋN�b��{�Ndl��:�e9tΨ�cn@G�q�{�g�R�����;��zl��g��48|)��0]#��Mı��ևS���L;����D���|>x�j��ph��F�83�~>��9�!��Éҁ�)����ÁD<���^V�� �QegLq�j �&,��V��\Ǐ3��&����۟�>wt;�*ꢪ�Px��96�)ꨇ%��6��|,�e"θ*��vX�oW����wX�4�X�)x�%|�n����*LJ��q��hǺ���>-������ �?�a�.�-g���Al�|�����kc�&);���[�Ќ�-�`�͔�Ĳ�YG|�ԯ�TA4=na�2v�@N����!�
���l�Q��_%����qMC�Ĵ2]�;���vo��T��xG����P�c��격�F��Dh$;sn�3��\s�-�5��%Y 3A�f�ɀ�'�ɗ�Yږ}�������d��0�`I�B��'Pϖ�5@�(1ք���t'���B�-2�-zx�&l�j�l k���ׅ��HB{?���P�O��Ѯ������
B��$�c��B@5����(��+�F��P��C�a%� Am~�Nbd���4��~� ���8��~ށ���s��P7Ѕ�Hx��7�d���#��W	S������Q"c3�혐��\�#�j�:��z	�n;����2,�S��0S�S?\�~{�cmB"�&]��ʯȻ@n�D�VD�1ݻʜ[:7��T~�5�]�+��VS�H�r��uA*��z˷��^�ꆆ��d��5�:Ӳ4/v6�oe��M�a��Ua�=�4ik;���v��6�=�vefhD�O�ݿ-)���K��&�Y�TL��$���q��1!�ܙ�~��:���>�h�9m�B�0��)h������ܸ�;O�����f,����Ӂ�=�U�����`B���JɉM�vB�������u�9}��7�a��G!, ���M�{3|%q!��jk��B����x�Q�  e�@k���M�����,7���?4�ϰ��Z���=3S]
���\߹93 �#(Mh�8?É|��P_�Ʊ�Qm���������aS����B*����2(��i��DE�������(�m+��Nj�AҤOX�p��p`�)���'��^��D,���E�e��u����W��k�pU���X�p��g?q&>o�	Q��՝3�x7����8H��3IkAR����t��d��-�Df�V�X�$ͣL�8���a� L��R�^�W�	�ڿ%�	w�3��ǿ�q��4��\����_|+b�~d>G�0�6�X�������ÔI�ǒ�Op�UEt��$�����Iv�.$���U;�����0�S���h�s��C�Гb��$�
��#����zv'�������
E2t�;pz ��) )/2+Ðvxo"����T�r��V�F�̩�4�nv
t4�����'��x���~����h���!V��|��G�s� ��Z�Im�핅P4+}.��g�����u0l���:c�ߔ�&P�{%~u�������Y�j�l�y`Dk0�1>Jk����M'G�k���V���ީ�/�=�v�%N$���)��@0���Q�X��"��\�KC%y�|�k��6̕���I\�R�*&vЋdS� �}>^�&�x*»LR},h"�S����̩����H��I��z����siH��;��?��!��e>]}��F�~��n��iQoϪ˨���zN�G��|��݂��h���$A��/U��aҗ	����˞��F��Z����NS1i~�'ԏ��#�F��$HUIS�T����PK   *��X�����   �!  /   images/4b131f3d-bb43-41b7-a007-3fb3641e8d39.pngmyg@SM�v�&(��EE@B�*�(��ޫ�ޤ�h#M:�""��  ���^����N�?�������svgg�yfvgO4L[����USU��.��GW(�����#w�jAA�
��S[
�M�j���I�KӎlA �5E�AP��T�;����ʆ�#8�x%�A�w�Q���6�r�+/��K�^)�C#����¸T͠ד���|�3�<,��,N!K�CW�'����ǣ#��v���-�嬆J�X攬����6ϭ�n�~N�-'�"N�T���c_0��	����|�����E���}�{lW�P�e���Ѥj��K�x�mĭ۷���t��7�}��(�#����� �!\58�8u�/��'.�L8�X�O��
r�g���,�C�!?���t�(���͉@^�7v���xA�(]��l,0ɰ�d�ge�b<\�$V'p\�������Ok(������[��4^I��G��|p�n����g��UV2�3a�8��DD
�J�M�?dt����N�%�L����j�(5�QM�>^��\T'�����&-�b!�MR�j}��^��Sc#��t	?�	�d����t8Y�^Ⓦw�B�ݭ<lְ�30}@��\���>~ʘ��Ӊs�CNT�K���>�y�^v�����Mb�0K�
�&���|�j��s��9<h��"/Z\�dOs���Z=�FҴ>���iV��
k̍�˝�b���Ff�䜅�TX����P��:ϫ}p7�����Ժ�<A^�i�@�/A��HՓ�"�������� ����q���]�QS�w����Ȍ�	�/�[�3�״�����a͹`3�$W�ayP��i�vwL?�d�����R�e]�Zʻ�v�⩍�7�_�G�G-N�c~9�6KYpD��U�4�_�]��g�+��.�D�,6��Ȩ���'yE�<%�"4���_��/h�-;��:v��ctR^��cUJ8��tBc)�� �Y�h�dǙ8���`{�Q/���se�c��~�a���B#��=����x-����$��Evz���j���S��@Ye?'T0��>cd}�s�dl�c� �e3MC�h�v?'�\��)&-m~�\�&�eģA&�i(��RG-a���_քck�(I�^
���4,��@�XǾ��O�oia�-	�zy�����*%S"�mn�&Z^��+���H�v���`'W��|��0AG�܇����#�2|r��K�.9�����Xp����'��դ��ז��>WL��B��Z����z�w�>�����-�u.�6�`KT��\�-(<*2��r�����5q�vR����pxd8�#=?T�`�c��'R�K��՚#�(�=z�%HjĚQ�J�cV��ޅ1{z�GIԓ-�*��zx;\K9S�ZE&4ť	�m���#R��o����^߈㓧�W'����uА��+R��v]D�w��[�@���^��[�%!��W���DKK{?E���V
J�eq �ah"6 D���)�j�ܖyK��Oܺ��Z�`F���&O$�W���a7]i��o��VVF'aV? �1H�N���8<�GoD�S����T�ƙ���]���k�|Nzf�}��|��1?j$�C>�æ�����mwt`�2y���3���۳�����m'l�����?M��v�Za][A�s�N����d<��<?/��C�{�&fdm�����	������5��>�L6�l��=���rR�'�9��sS��'���h(&8�8�r�V���1Ԝ��&���:��Ǔk��IGc���0+B���z_2����MR�	n�AZ|h����e+Q��V��P@@ �� N������F�4�����:G��<�?;;�ܺu��+**jdyc��tg�b�s�t��b)y�r�/ԛ)]l� `�-��p�~��4���W(�P=��B&���W��>q�9({
���joy���,%�3_>^�dV��;��8�'�K���gQA����єo�r��T��jU���k{G#�Z��C#5����͇u�eؖ�+��o�T��v)�_l@:�}ɣ���v�_xBe~��(-%����4�&&'W`���с}M�v�BGQ��UD���i�S�sLIjj��U����k�Z뿠W嫟䠁�k��OKO�Q����l�,�]e<F�n[{��0�}u7���W�#1}���yx=DBJ����<�d�&V�,������-p�g+�xvk�k�'��ƫ�:!�{� �+��;EОԄ�P�����^����~hqS�� � ���'�C�S�'�4�~hWsQ���j��#���#�����˾)F<���j:�u�*>r�8����7T���/36�T]kC�SW��{���AS^*��ή��Lp�� c�2��zJq�-mC�צý���s�jw~�������R�u��W2�(�%�l��--�qE[M��q	;c}�Q<��T����{À���v,Ș�ۖ�0mE65�h�"c.�n����%�|�v~8Y�w�^Iׄ��F?3bv��j��OPv��݋�͒�����P^۳gLw���4��qק�YY����[#T��������=���;:��JT�ɥ@��Iu-��D�]��7$mے[�t޲'Ӳ��oa�P���,��|��>�F|�� ��;{���<Ԫ��L��̂�4T�@�/0��ZJ�T�j��˚��Uq��f��2�=�D8d6�yx7��{ݨ-���W�:"��N�r1��INVH��*���%s���en^{U9�����u�����
�G��<ߚ,�M�R��S(�!�3�6��u�7�ߑ�Ui�='6J3K��Gko�?kXI�m1��	3����m�{%%i��nw��Q�Bx�QKj[+��4O1��N7��-��b���	)#/�^��#�%�r6�:64�rs���}�95k��/�Z�Ԥ��wf�dJ�\\�ƚ5��5T!1_95�=Bוeu( C�[a,��&�F���ɽX/g�Ҹ���*$��
e��rCbg K��+E���uڦ�����4`�]������jz�zU�vZ�YKY�c���U��o�z6�Z>� �v��+++L
�g����ɕ5�<^�
}$W48"�Jt�V�P�4�L��0��~�~�}�̪��Z�c6݊� �� ���͡��|ھ���Px��X�b��V�H�F!L����b��G����ngy��M�{{��O䀝�_jZ�^Y��6-=J�<�xfMXf��`��5�-苼�i�߿��H�/!+��H��V�6g�q����?���6�z��5w��WG�[Ͱƣ�M)�^�%�s�#1�	�ݦ�E��=h��U�m.( 箋)58ѕ�]ӽ�H���sd��=ճ�6s��Sd��{j�7��Oi�k�i��?����yR���qL	F�<
*2�	��0ٲ�'ڂ&{J�<�@ �X. I��@
��%|��^�v�RsOG=��s�@RTG.�����۳l_��nt_@D׷��a��=)%,d$�E,�SS����V;iƺ�M�|	K����e�����=n����j��!&�ݮ���A���ͷ�-u|_�I������R���Nj�C�ޥW�e��`8��8�HF[9z����i���[���@�<7��lj�f2�r��#�����`�+B梯��������:�ϊ�y���OB����:� �B�g�_��^�f�z�̓Lʦ�o1��ucc� �VC��.�*��r����𘏑�SR�t[m0��J���S��m����|:u�2��E���	�o�8oM:����t-T5�Xe�b��Q���Qt����~:��=}pS$�?�ꑾ�he�T~�&h�w����������?M��]7���֑'�si��Gp`K{��x�I�����BTW�Sp}�Ø讕��eJ`��zժE�L��GG��D�v��l�[�LY���8�V�����K.�[D)�l=�5�.�c���^�Α�s�����~��lj�z�`��E@L����g��oN˖�`�m�����[0����r��d�� ��D�f�Xe�
z�۵gU��G�!d��w=�����2\2��y�f0�&�/�̥�\�W���E��W�[h�1|@Ǵ��D��G��<�OH3S��?��̖4�VL��9T�@�ͮ|�E�}����}<����`�'�2�͒d�.e�=�m��"W��2
,f_cb�}�h�ε��G���n �	����q�I'��-������‭F�wL%��f�=�	`bC���^F�Tf��!�LO�,�j��puqQ���+���@����>�n1��'�O�\Q� �;��c�L����I�Q2�߸��6z�c�Ziǂ�
��|�kM���zkZ<Zt�od!�N��T�LKQY�Aw1����ӽ��	�
W���g�ڽ���V����h:�CtH�����P���W;�AS�ΐ�Ō7�]�pI���5$��YyLT[��rrR7D6�f��A�~>�do�i<��`C��5u���>�kA'��>:�4��*����m {���τ�N�X�<��a��9�S���S���[@�p��HyR�?�3�AO�U���}��k����2a��g�R�g�q>�z+�{I	�S��F���e��a;�ء!e�r����ꃒ3	-�ځ�gV��gc�2�Y!�j�[;��R�d�� �J�:�cT�S�Uz���G�����-�u!��	̋0'�Ѕ8�Ȟ���g���7��2A<�_�K�F�^������ކA�#<?+h�E�6�ج��ĸ��Q߬����l;H�f�t�T6"c%�ܰ�>�f��N�s�.5B.�m� Mi+4�u��@��`,�;����Ճ�e�g�G�o�'*J�ݑ�U�=�<��?��Z�	j�$��os����F-.A���J���/�;ܺ}$���t���A��6uL��pn�����i�b�w�C�]�o�E���: ��!Ic(K"��~Z^g�'J}��#o����""!Q���;]�ٳ~�֥���w�hٔ׭i��3|�0�[
���g��Myi��Bx����/M}�-����&%�s�F`Dm���M�l�k�٫�g���$w���犂�dl�Zū|���c����J�z�����W�I0ԗ�lW�̡¾sHRˡ�gD%{���ყ��KjZ��A}Mh�y�6�m�*��G݊��>�&[�x�.���V5ǆ���ӞgYƬ~n��þ����@��ЀQ#?)Q���W������?�C�*w��+>"��iT[��&r�$��q�k쵷���>XmR���-&s�����H��j���GBg!�S	+G*.ldK�P刏1��N���\k�Ā���<�AhI�|����QGW���gr�Jv�@a{��Mv���I!NLӫ �|�
q��W��^�ݭ�b����Fݥ5-h��_E݆AO�E)�S�q.OR��a�wC.H��L�0@�LF�h	����#ԹX���ܩ�7�7�+�kשZ�[��z����)���U��߯�@�euypnU�4F@r�c�:�q
	b���&V�$��_�j�-^�Z�P�k��}�ǆ�JU҂��y|��1�t̪Kau��dJLLT�v���Xh����s06t��z�u�|i�ALȾ������YC�u��?1���m�2y��*�<Wf��1![���>f��I)���Wnh�o���s����s��(3�'�0ClD{���0�Aj_�z1#�S�5��9��b�>=��{��v�-淉�}�ݻ�z�/�Y-����ӟ.�Rm���ә:'���;����'�5����>������m&�ʼ���0�̐����l�|
 ��Kr.�f��ؘ���﷧�,�!{��f�*,����k#�wA>d�;i?�S�o�������j�+�|�h.�S\1#\�Z�>:���[�}^�p�P�^�B�w96t\aqX���8��iKLC����΅�?紣�����{y(�seű�����󛣂�G1UmB��G�?���̚���=�')�EfW'Vm-�5�T`��
Y="�nii��k����b��\��5݉�*l{Qӄ����41���q��Ϡ6���[ob[�b[o��ZUz<s��_��樏a�,t�y{t��q��5��Qii�?�V��y�Fk��l�N����ni���f	C���1TA-}UK��7�h��8q��9����i���'xLD"�GަO�
�6oJ�k�L� Jz3$K>�]��%�E�V�l��8D[�9W�5y����-�u�u��+����p�����b�}����͝�R顂�ۦg�����K��K�T�\���7� ��g�p��1�#*����4�3�.��x�3�_�DD��򓭦��W��*n����#��M;_ƿ��U9t�f����9T-���>Xt�����E�sq�ݭڄ��7!&f8���bn(}�#���M1�g���L��O�t�ſ�]6�r�X������(��o��?v�X�n���/c?��.d�<E���Ƨw~�g:B}�������ܖ!kn�0d��,���0�.��@��esN��uF�����PͿ[���;W��%�/R-v��˽_�?<~����{$^��-����������6i��D�W����a�T�~�C��c��1���m���~5�6�_�o�͚� t�F��1bQi���y���>�N<:U��hxOǛΈ쵑H3�f�ٓ��gXGUa+o���)+�e�=D�_�ws~�(���ȇͭ^���!����M��>����Q!N������ �"�*����F�sl���y�Zvԯ��W1�nR�d�_)��6� �Mu��WyJ�Փ[]\K��I�Ei��f	Oa�L^}�3�y�l�Ĕ}I��Ѽ�E�ʬtx����?��;H����^~i��Z]���=�H5ʏZ�E|��(����T{�֑�[��!��
���VH�1�
7���� ڤ́��;^%��6�/f����|<�iuZ=^[XE��>V�ɍ�"݀��7��EwIb�1mO�����K h����:�5i��9^�E�:���߀�x4�m@�9����tL#H��f����~#�$�w��t�suph_�2گ1�I�c]��\L$ �5k�N�A�f 3"��sH�dpR�W�^h5�H�$�����������*�v;kv'`r:�����c��$abH�2-�x��x�"M�|>I�h_wÀ�G�q���E6��h5���v�����w/�������xRhp�$�����I���WVV���fw S;:;˥�����EZ2݂�"���RgL[忟.�Iz+�9�aL3��H�Њp�,�;��ɯw���O@��߆��9��NX��r��7zE>a�'K��b����:8+.abL*"$��k�^�E�W�/�<�&�zʀ��=֒!X/��c�'��rIgU�u��\���������$���Թ�Hl�Cs.:��D1h� `���x�PN���׆�����SQ��
�%��t��t1����7�z��v;廁��bL��R)�P�Mzdp؟�oS��EwG^�]��}���D.�C��R��G�=R�z�T#�)���iy{�L���1���Ec ���L���$�M�F�*XQ�%�Q���@W�Тq�jCx�t�I�"�P��\�$�?*���z2�#I��B]��E��t�%�t
����D~��h�8�Ӏ�E(��)�d�2�0UA��ܙR%W@/��хCC���0�C��dL�]��'Z��DF�R�(��-
���"�1�> е[@9���	�%E��N*�:�T��O���o�*����Ƀ��J�i��Ѫ?
Hv1�#<�C~Z�q��
�_��@
���r�G��NH��
��$�H&QXI'�|��l���M�!J��������@�j������V���_~��&7�\h��FO�#��Ph~+{�<FT(X���`�6��y�p K�s.�l��u�>��W}�\0����g�	�!y#�֍����z�u���@q�1r.�'G����K ><��T�U���#�!�-PT���n7g?!-�G�+z<�����m��[�L��G;�qsuN�8:��TW��\�,r�2c�"�F���5��˖�Ӑ��O�>n�r��%��t�K;�כ�:/��eh�<6/�^yIz���	��+�HY��¤@���΍K �.����R�A+C��4�+E^d\ɋ@�+��u����,Ћ|T�$e��;$6��S����j)#^u=�"���NE��O�`���+�nM�zT�I]<�)i+~}b��PK   *��Xj���(  *  /   images/6c8b06c1-8935-4e1c-b7d7-4989f9141afd.pngm�uXTm�7:*�c�� �"C�  H�H7H��0Ð"��C��RC��tww�PC}{����s�?��{Ͻ׽z���A����<���K}x�]g��n�V^J�w�IY����z�!0���������4�@ g�ߵ)S:w��@꽨�;ts�#�Z����]'�����(1f���p�'����σ내�ߚ>��	����jy��q��l�$R�Zj]S��x��c�J��_ٚ�����ht5m��^�\:ݭ���ȳl�U98,`+v23+�ϗ��zNb?�l�#����-A��I��B�S�j׀	��;��rrr��������Y_�~�������Z��7����4-��~�9&��˽�y��9.�5SVV���k`�"��ں�dr,��VFKK�|�?�F�P�l
lm�D���l:&zwסb���ka��aa����VbRRR��IN���[t�؊ҡ����cWed�S6�-{{��8.�鞎�������VXH_b�kx�+M"�#M��?�5�C����^[M����)ZZ��G��%|QUuo�@LL��&�,�V!��Str�W���F9�:� ��:��֯�Y�^as��Ȍ�t�j=���6adZm�2���)��~c?qR��Ü�ʓ��n��9]|�/�rz���t��g������j���\:vB2`C,�����1D�N�p{d�5�C��Y/*�־�M��k>�ܢ�uW�ջr���҅�bҜ��� 5AXp����g��*�C`�x<��e�QbE{��T��`����{X�$F�
cTZ���)=��31���S��g|Kb�:PX��7L�c�t���d�#��?�@C���O-��MO�$��0�� ����	�7��m'���'LYt���F�(�,������/{g����`�m�����*�[c�%������2��b5�-J�\���z� F����>������'jĉ�#ba�|�;�=M���\9.�vt]9�k�!���Jm%�3�}����N���;�<�[ZY�������M�����Q�������uS%jy�goɣ�Ǡp����1m5T���^�ŵ��T�q96'0b*������J�SK@�u���O�~=���´��ziq)�F�Ģ���XL�,�����e������Y�^)�0���/=�=�7�+N�(~�O�L�H?{tt�ڨ�6������F���0mH�M1평mt{����Vz�������7��_r�2���!�R���"[M܏��|��lHθ'����xΔ�/��'��d�el�h�EE�靟�u�k��'^����+Oп��m����p��XX|z*� �b7Y����E�P!u�����,���Ó�,�EF��z�g�\�����n�h2�R�i���hk�b<��.��R�s��r2�x O|�؄A�E��H���<�>TEP<�Jc����������Ư�1w5`�[%?�j���ܺUc�h�����΃�:�XϜH,I�$�v�w*��`Y�tP���K��)�+* �:�H)�1���f!�J�����K�!��?����%5wT�Zrc9��)�NH�7�5ʰ4r��~F�K����X[w��J�}@JяJcI�������ʵ'^	�2T��pv��Or��ĝ��+�̜r�1�$�ldo���85t�q�Qל0��8c�99�0��#�Sŝ��{�7i�<gu��E�6��{G��!�9�/�<�C��9,,IvC�I<���ϝ��{J�g�h|R�
ޗm3I�����䟂��G ��(Lȇ�_��f�"�zz�I�.��)�O�m��-�Dt[�l�;3�F16� �g�J����nCӺvB®?���n������9
��������^t�9�9
�C��癜��5KM�򡵪ZZ�Z�;K���^�|d�_֐12
@��/�'ˣ�W���Tωh7�R�74�>��҆L_V�,��(��*���Ƕ�Y��e)���(C�O�R� ��
9Mj�X Qk09kf��Kg����u�]�QSާM�����MX�ْ5hԞ9�NpbV�wb�^��.ˎs�$���"�Z�%����}������ivZڵ#M5�[9Խ�͵���A�>�:_��q"F���{4]�[�V���?���B�;�Mu[��\�X.��r�ӗ�gY��*B�_���E���q/�����΀V�םt�I[YY�d��)K��K}k�6PD�)�qo�9o$��5�7�E|���tQ��#����(�,��c���2C�N-\3��(���{'�U���0�	�6��(.�qldۘ��>oy���4{��"����ʓ�V�d�SZSR*~)�Ɂ</-�(����ujPkؒ�8�0�4�s-W?F�w^�^'.<��U����)������[s����ʆUא��JNn�<��y�y�VH�ňU�76�G���� L���W��#u~��	�~��,������58J�搬^��Hz����<vXc�钣��Ҵ�u��ÚW�������.ѥ��UT�V#�

�~�lf�a23�����P����E�
�p�����g�g�7�k�g�1[tU�l1�_u6��ʍ�����j9Wc����\{l{��xzN�q��Vl��H�H&�>[�v�ه��;�s��1._��@[8iݰ�Eo9��5ic��#�a'm[�7�>B��^�2O��M�p�Ō�s���w�$||�cL��ΜⱿT�$�^Z�Xeܪ�y�^�!���3�axh�C�_핆k�������tl�K��]�W�>��1H.��w�4=���Q��:]���-�'�G��0W����K��]�*TH+:+s]�|GnO��f�ĝ��_�k��v��>l!�9����/��h<�&{�q�ynp�okbՍ�m���꛻)��Y8_1}�K�*��uyR?�]�[d=����Y�U�vRs�K2͜�$:`�[������1�Q��#��㲯_��F���n�������3DapQ���mcA�q�N9룿ce�oݝ3Ղ_�NM�|]�QJ�(�yq!�|W���yO�Ta=*�Y���%�4�AL"��
)~���o`���8N�����P���C��2\h�y�E߈mM�������� Nٳ���m)�`��k�ġ�!�qvڍ��܎�퐮�~�u�!�sIŢ�}(:��������<6�}�!�9�ʩ
�\1'U������E�w��p4�썖.cL ���$~��|���^���I5����.�ޏB�\�kH%�M1<bҔaf�qq����-^�z�ǀ���H�9��k-�!�]+�D�����2��y���	���a���A �Y	'�Кe���\3�� 	��!�cg�*���L�7�l,ۉț��d�Ԙ����j_�IHN���;��i�o�H��T}���z�C�NTr�T|�;�+f}9����H�3�%�.dYw�]o_�v�_$����p}�x��׍*����c�"�#G�3�x̨�5(���M�I:ò敝7���w��l��,KM��wz��s\����4�����t��]a��:�a��84va�� ;�_Hd�m �b1�Ly+{�;���|�CM;�DG��qv_�������&
��?s�I�����OR�A��ۺ���6�-8A��}�vu��@X^w�d#V 6��̣���5�	]�Aڶ'%QHYʻA�cv�u��������>�����gw�.ͨ����N���L�"-ǽ����\��)paF�0�����4 h�W�RO~Q�3i@=2�#m��?��D|��[x(-'W�W�f�'�#/-M��-\R���ϟ�2j湅C��&������,�L��f¯c�|���[wv��fb�~��J}9��[����[��y:�b_TX�r?]�7T��:�'7����!��W���z{,S�f�w����c;�~���"��6(�����[��Eٛ�}[�L�6��\e@PV���m!���^$�f��J�ۣu��zT����K_S椚�U##4�_y�̱1Z{���G��{��?z�`;���AO~�Fm�B���@?�֦�A�:�+X��k��=4�%x�~�X���Cm��޳N����y����ܼ>��1�5��e��\���@��Ġ���Թ�>�\L�*���=�0��g��@O���#"� .n�� 2�5$�{�0�B����D丁K꜡/+�����U�G%ITv�Q؃P)����x�2���yb3������{Y	��ze�߷�S֠�X�	P8g4eg�S�+V�Fa��e45�	@�^�BDj��$7(�+o�>���@$�����ZC�tmP��LQ�IA@S�e��"�x��Ҭ�E�����e�o;��h��r;���/��3��cJ""�o|j sR�Y���Y��:呅5�&���q�l��{[���b�8��m+bm�xᮡ�D����Z��Z�d��KJyE��6%@	�~z���6����T78��GPO���(��)�SU�I\\\��n�v�y�C��,� ���$�"E��uעu�,���PV��9:放�4���$����O�-ϭa*m�S>���5��W1��`'o�7�� 2�*Q��N$�&,��"I�^x�*�C���E�{Et�!}��#[��<+��h�jk�����HF�ܺ%������v+���%]dP��Y�cJ�@��W��r���,�ve��]ğө����y\@������hmm�B�v����ڡ�5�����1�њ��ĘA�B�pN��A�����)���n�>��R5��N�2qq/��"�}� �ΐ�/�o{���h17���?]w��2Y�?�Ғ���-��f��?�hO���J�/�}�a~��Ѹ �ʲ���6����}�6G[DU;���}ll^V�K�&�&�#K�v�p��=�ڄ���򂂂J�";��mDʌ�s��rg4�l��jHZ��K��0kZf�7:�{��nn�x,ҝ�_b=�)�N4%��am���(�W�}�;E���պ�o�?�ID��Oև��N���� LU��'����k��#��+e�����n�Y�؈`���d-�"��~{�{���q��Q�tÊ�l_�?��E!;�<��\Q����%B������= ~edg�!W2n�y��P<�H�sQm��:���@��-�I��YEp����mQ�ăE2��-�"Wh����:�����FB�~�� =I�{,��w˸���l?��m��:b2\3f�j�(3��(����`�/"�!PFǂZ}==3�)�H,6)2;�b�`U�͟~����+��
�=�ء��J����2���.�2( 8¼�H�������'y_�h��
j�i4Nؚ�1�T������ʍ��͊.[###yyEf��C��ʎ��gam��2�e9H���?7�vvٌ"�;K�GL�>3��w�~ռY׽�y��].�y-g�a��ʏj갱�,_��۪�=V�G�g��O+&]s���V�7�Y�M:ᓺ�{���#�2����q��u�6**օ��k��a!��?��F+��ݶ�g�M)��݈��C����#X�wzKA+��ړ�i�G��چP��!:/	�z�F4O��Z���V����Ym~a��h�v��ꆆFܷ��ɔ�ʏ1H�"���M�"��iNx�O�=ln��t��z�u<�dD��z���q�;��� I<ܽ��_OdQ�_�}��\n�+<(/7q�B�L:��al�j675��c�fqgs�-���˅"��矝��\Z �a����8�ⵗ�r�/��K�ui,���D�	TN���_t� 4.���儷zW����_Vי�+��N�\���Y|��jC���89��˞��m*�?^�*��S��$�m�	��e��q�8��l2LՂ�30�9qj���]�u�g�z���u$���ƢI3T}C	`���~�мO�-�[zz���Nȳh���u��&��D��88��"���l�I��<O����6k8�T&�2�6��Vt`h:t�w�./bj��1��(8;�ꁾ�}���Q�х�8��p]��_$�BV5����\�!!I��"N>�r�Mi�����Ŷ���~w[;:G>�Vh�����Igؾo��;כ�K��B�4��rC<�=��0\���m�_�����G����ϡv�V)L/{�k�u˅v�u^��-[��*� BB�!�����S����ݜꗯ�j��P�4�(��W^G���oj�[ם-��>��)}�H�"=��s�֭=�'B<
�bX��z<�9�q�N���#|@,D�y,���˛E�ָ���zsm.�s�M+G��J\�'��o8�=%���Z��S�=R����yb8:Io�߿�Ƕm ��_[�ow`��%���{�H>yh��;�ݚͭyX��ɪ3��k�^W�~�}��II�D:em.!O��p��>�b?NF�#>Z@��[���]i?{j��hF=���[ټu�������i�E�-�S0Q�q#3?u�q�-\���]�c��ӱ驗�Yk7��	����D�!L	�k��Jl�h���y�JIG�2����{3�KJ�Nn�X�ܳ���ly���4���	{� �%J/��?)qo��b��}�S[��ڒg�׻ ��r+����۞��'�ԋ�S͗ė��K�m���46�8�6i�٣iE.��ů��tn���yE����'��FHXC:�l��CCM�{�}OI_9���$��9!�q(w�ꊻ��{�\���-o���Q
=*��ALb�]ڊ
�/B�_TO����+��v���l���b&��w�u���Lܼ��W�Wag�q[NpN���i���V��A��X{X�r���G�s�thO�'��j?A��dJ�X�_f5l�c�Q��2zq�^'�n��66｛'#��ڶ��ν�vLl���v��{�'.)�%��߭�*����>��([�,_5�{�nD#���V%��tN�=k��ŜM[;�<qG�[�b8�-;��sD�[�b_���2�'�P٥Z����m��\�W,���{ֶz	?����,��]��_/��
��b�y���uߟL�L�K'�zGABl��ߊ~I�E���ь��S�&��W���8��*B�Ul��V���M$S ;��R)�>K����q�V�U>��ü���7o�=O��ygU�%�;|*�k_pd:�%W�@SòLFj������
Y���~��/�$a�+�}*�{6b0(t&�EL�i=�^�1.<B�����\�C�t�*�BM_e�[����@��4Avv�L�[碊���{i*Y�T�{��h~[�
�D�ݕf�������Ҩ���D�h߂��F Ovp�����sy���
�u�>�g�aa��-er"��"uj�g-��N��wɈ��޻�
���2h�e�߳v�� R���T��N(��}�ml�[z�[����y��QrE[����Ӛ��\�m��M��c��n��h�ʪX$l׾��j$;y�Z��tPI;�W.bSR&�H�����t"����S!	��mg�z�.[�1lV�%��j�{��U숎�o)V�%3L9�r�n�i�����BWT��ky;��s~�MN8�
��N"���ýϾ��y�5]��fFUlY���)Ș-[9�`(TG硧�6��J$'���Kၿ
����ذ������űu;��ݍ#��Ե:
˴������h5���K������m�XD��\/b��h�=7��c+M�r��"��NB��w`=�t^SN[���~�v�|!a}�-q�9WO!��s>��>����yH�R�Sԏ��O6�l���C�՛V)�4	ĤSz�+y �Qɛ;��h���y�y�]�}*�~���܊i��-�(̐~y�SQ�ӿ�R�x# ����i#㠞z�<��A�S�I�]Ϸ�oM�d���дtp�S��,�S�U���{Vk��r�a�>�Ps���v6��5����F����o�M���+����E����0]�)�\�lQE�ΔR5�kw�a��Ǻmk}l�|�ڭPu����d����)���V��	ŵ���w�rLt��j	/v�͖�d
�P�#�c�g�aԇ-�w�l^;�2g�W�<v��Yy�H{���JC��ɬ�Y�-�k(��)	���苊i3(� 塖���1��,�\�~�do�ۋ���� �[�&չ4H����x0��{�D"'i6�Bi��tF�5T˧n��u��{u�:롤���D�g���XV]�R��ա�r�߉���'|�ŕ^z/V�t����LMo,���v
wmau�?�8	��=r3���٧G�5��hD�샑`���f�����G9��+e-+?bV�i�@��ޮ�gDJ�I�4˲u�*��AHH�`tӹ'����yͧjX�\,�.��?J.�:�*��GFt�i�৮UKcT�.�Z��?��E.C.���v�C��
(�`cd�&_#�3�.��M�e�Y�(<\��h�Ő+}�vW��xCx;$9�S��#?�D�f��{�a�J�֓�����~�{"�G|��gZ��gPO��Sb�XZE%+IX��?8T.ۥ�VP�եo�E���ձi(��{��c!�Ƌ�T:��;;k0zL�����j�y��w�=�=���B��1�7!8���;j_9��������.��A�a��A� >�z�b�C���-׷`j,��@��<̥o���}�ϣozz��l:��5+����,��Ay�gK��=�{h���?}"c��:���k"Ŷ�w^N���vy�5W�=�k���?ٻ�^�;��)n�r�Q$ 9�H���<P�:��u/}ѵ���`ijI��g���^�ُ'���:���>Y���%�3=5��kT����������Nk3�A E�s��$ �����[�@>U�hqT"r�֢0pp)ԡ��6h������حs�`z�q�i�	 ��e���!<�>(�@o#j���*E��Q_�H��%� zP~#3-������.�(��>~c������k�������^��4"NJ�zRy��1�8Q���j�~�yu��
�(!)9	P{��Y�54��̽,=^
�sX��u�G pUUՑ^�w~���M�Y2@Ew� _ϟ��u���^�t�VH�s�s(��)����3��GWn�����Ϗ :����E�gȈ)Z�?�\В�~��b8s�!�^)�+���W�Q���95����Jzz��Gܒ�\!%�w��.�7q��1�=KKnQ�C�]{��?�� T�,�w�4{O�ɨ�IqE��9e�x���J/���I�6{�3�^�C�]�nѧ�m)m�Wj5�J�cB$�/�.�{��]W�e>��.��,,,���m��e2b�����E��ػ�*�-^}��'�%�-�qjx�2��K&��I�#ݦ�������{�t�}���å��+	W�@^��RҖ/?&�Gl
�9e֠O���Р5:$?Wr_��@ gZ��d�\�]>C��W�s���&�C������^����1r�h1�0�m0�JT
��F{���^������Z�R����i��Xs���*��*�\�h��;^3�a�%0�o)��
�<�����v�� ��9@���" ��HK��'98���(^�;���/ ss�%^"y�����y?�=���/зLFf�R��GKI0��ҝM�N~���)�?K�m�\�Β)|RH~J�J�"4TN�\��
0�
�L�U��}�;�)E��+Ek�=5�����)V%��d,�G��5�&�qCq���L��Y��f%����i��/�n��Gyf��ڜHM�Z����T���^�@���2po��J���BLAjy��h��}O�s��H�hY�8bC����`�BNZ9��#��z�@bu�{H�J�؞h�Ft5���9����M�l����>���$_�Џ6g{�s;�?NF�L$Iz�4�, p~"��F�U�R\��H�Y��p�Q������������HluE���|\:v��-\�� A�ႁG%(+)E�k�#��E-��Ec��f+@��:�P<��o��B�y����,�ʘ� ot��C��%�TA0�<M�\4��,�?�~��D���\�6��J��{Q%�cٰ��6���b��>�6����xB8�cl�W�`4>����q|��߄���u���bN��:Q-F�q�05�������
�&�EDx��q��ݡ4��Gڽr���-r�؂�����.�J�����#��o�>��Q�W	8�����{�׈JG
��>@R�������PK   |��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   |��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   |��X#�@�9� �( /   images/bb1d7dd6-69b0-4e8d-a72d-bbaa9fc3070c.png�eT�m�7:��� %��1��t�twH��t�" �t
H���"u"%�Cw
C���<���{��q�^�B/�9��<�w�y��&����� ��ܘ�@��o�;��R�pݥu���?����-Cw����a��nއ������^�nV///.['{ws+.g7��m�-DQ橎w��O�#��{y��	^�����}.ߡM� �ħO���g�M5�ޢ������`ʝO������S)C&�J�Y�D�MCc�6݃�䞿p��i��A����m_:E}�Z,Ho�F��B!�g�!�W��ʐP%��y}�3�G���k��v��I4���f��뿷ŤP���ƃMa��z"��%ԙ.x��l��?����_��,���9���mN?�,�#g�ߚ�D��ʀj���� wm��ߡ�?L��s�{�+ބ���}o�-�L�4'�;mY��iD��o�q ��Z:o�)y��G6&�i-P��~B뜰(��/m�a#���h�h��!�:�6'�~��Ja[�.��0�ū��|���1������.��=��� �r[ f;�VW�GI���r(���1'e�G�
�6a�@wq��)�{�uc��Z5ʿ�k�g���$�Dx�{�e{�H寞�8��J����3m�U�P8m>&+�{b�~��"h��T<�s@ �X��q8�Ѕ=�XxxW.�⤊Ʉ���S�}�Љ�4ߊ��R�7�1}l�y�ͣ��5g�U�,� �'M39j�X�+�T*t� -�#���KB5F���\9�Ϳ�=��q��6��:(.���<	�&����/~���
ўF�\b������L��NTvw�%�h-
`lE͜�"R�� ���	�zS�����u�rL�����v�ʟ��r�1������	�����_�OKZ��-����D���om9rX��Ĳ=v��K�434TQ� �'����(Qa�J��ܵ������_{)W��V���=Lxҁҭq��0���5a$+��]�0pȵ28�쳮���t8��cbb2;5�mt�\y¡�f(K֙�(�D�y�6E�A�i���q%����^^��}�&��/}�G6���T�	ŝZ��G�*G�9���F��Cvy������u�Ү�<Ĩ�!;�Q$}��^^;�����>e�ͥ�\^^4�۷�v�1x���B ��O�l��t��d�F��=�ä ���l`5F�*5� �?X�!��G��r�.�
0̜s�*�Coa�q�mA �4��{6�`�)h_�K���a�C�l(!��m�|95й�{@���y�}��a[�$�UsA�hc{��y>!W�FM�=v%1�?�F����$w�c�c:�H�mxr2��?�k����\�y{�!3R��V('Ä�bC��C������A 	[��~�M��܏�����p��:T�
��c�k�ba���1D�1���ȝ������װ.�x�8�2��c _����y͸����\"�M�z�G]�\�|Pp����m)��z@ޘ��⿨����Ç-OF�'k�Kkkk�?	<���<Ǝ7����7](��q-�b;��~c ��
�dg���K�;��$P�=�r��b.l�� �=�9�s��:��ׅ�����m_G�m�A��.6�ׁ�+��|q�ݦ/���W���P��n����m�ԝW�t1�&�Q���I�4��s��3i��0n$�:�L 큟�a��O�m�>��Oؗ�WnBn�מ������G��ֹV�54h�0�V���2�cAZY�%���i�3m �����o��P�v,�sHUv{�Q ���04�c�p�l�8.�(������
�*��H�}m��{B���$0����b�.!��	Ʊ`�4���+f�ؐ�-�y�4�K#�&��A聬��Y>����xY�W�3����aH�Ѕ4n}XI��I�p/^�e�Rt�tD��pE�U�6��9_GW}���/��IX��K��������/��=ML�o�B 5սk[���2�T���Vg1�ߖe=عR���j�Ɣ�����hxU����ӞtAw���RxE���(�3ߥ�6$_'��*^�o�gN+� �	������I��'$c(����k�I�o�I}�6�]��n�Rc����U�r�"���o���ђ��ēY��J��ã����1�����P�d����2߁��N"����<�(��Z)E�;>Ѷ;�A�+_�w8��*�g5v�T�
]_]�M�Rq�ĪK��IIMe��"Z�_I^-
����hR�hY������(U���J{��DT^=X�;b�� L���Ԃ�Į�{����Z���J�k�+ÙҘ�����r���2��0Jj'gf��<�i8Z]YhOa�����y�(�"��%/}��w*�R���+�x���~�t�-�S���AX�J�>m-	��^���_�L�S%�C�hM���� ��.�8����۵��S��/�gGп��}М�ѐ�k�cR�6E��y
Y�e1Y(5gQ�B�>��[�B�H�!*@�}��w �d�<*e/Ψ�.��u��'8���j���U�Ƃ�>*X͙D���U}�s�Ѵ3N݌�ۇ�{W#��^�${���׉�}���Y�(W�£��?�w�d²���Eg_�tW>�m�=�J��nl�A�����]�g���
/ߧ]PX���/��������V��Ҡ���5k��T:�]j�xl���+4=�g�~;Ql���h����x̊��9j��������q��U��=�_x�����_<�D9E�ce�v����㵤Z��P��&E�U���*�i'y��;��1���o�u��y��zx�����s�{,	!�Q1b6�@6�9�1E�0�r����.��)��XNBu������>{�_T���Ao�D��u�	����a� �Y��1>�w. 2�X}˚��И�^�BWĶ�K������bt@����fT��s���2i+����G���$������8�6LMj�;��{
w���s��H�X0)j�\��䰒�tX3�2�g�FV<�4�S�D�~�\�)H�׌�����8����M /�7A����&�)1Y�������)� GcÏ�`�hG/�-��TV\|3U��ް���2{�������g/s�L:���q����h1������gK���OV4�s�A8���؆H�R=��c����h�8I����J�vmrӽ��)29,W5O��)�]���8����O\#�>��"��O8�)'p�-�$$ԑ�c92>�g�a-B�["ٴ�N���,��3-b���DiQlw�0���Zá�"�m3]���閟	�ۯ�c�3O��>B�nܶ��8�w�+�49�P�F�� ��-����x`����B��'��(N��.�?���rj���x 9)����Θ-Y�L��s�:��Qt��KH��Y�{h�i\��XHBh�y~�<9=o)ݪ��?��Bd���\��	��F��-��Ԧ�~ͣרCs\���MV�od�u���^���G��gQ�nR�A�Z��tĐ�L<J"X/~rrp+Ξ��Sl�gQ倠 �i�,���+&b��a�x�V�`�x���R��6>Tw�_L���\�Ɵ�y1k]�=5��Z�L�	�q�W�����Ó��ʉv��D��<~ܷ�a� n���ԼI�FU���T����/z�K����G�1�>��+|�S_v�&YGF6{��t��W��/��*3a�z�z����򰜪��3��4�z����N��Ϡ	b"m�2�Y�E��~���E]���=��g�+R;�X��+��􄤯[1�z��|��[���r��+{��Ɲ��ʀ��\y]4A�+A��φ]!q�4��x&ި�f��qW�*�1��.�'O^��p�+qJ+5��Gu�Z��Lz��8�%^�C7��[%��#��ޝs���,��¹ C�˩Rb�逢?e-*��s����>�����4��s+�6���|�����]�aտ9Q�o����`՗�V��5\5(aO��7ܰ�`7�1�'�ӄNU�g5��~�7p"��oBk3�kNӱ���9<��3+�r"e�޸N?ç�rE�Εs �xّ}s��ƺy�=���G}���8LĊ����;8bj7t�뎋{�/,-�Ə��|^?�C��ǻ��<��T,Xt�O��K���怤��t�w��"�Y,Z��C �M|��}��WT�Y��H�k�%rBs75jHT=�9�M��%����rnF
P���}XF�
�y_���3yV���j�و �.t�E!Tn1�[{r����hh��C[3�وA_��AWE��Z����YW�	�R���?/)���H��g�5�{a#ڧ"^��g}���hO��E��D�U��_ʔ�r�]Xs�����_s~6͒��S˫�k����z����z���-�\� L��ϟ91���"*q���N����EediSs����H酡j	���G�e�%S��,}�KW������,9.��Zn&�}	0� D%�2��W�����$l�$:��0uj����j�[;��z=��UKC�gX��z6��L�Z�F�;�c��{UѬ�ߝ�}�k+�RN�n����.�.�iy�%�,��Q9MSX��G��~4���7l7l�����p(�zb�N�j[JF��c�:�){���zr�6&�� 6�HFN����L�����[Z�ȸ��꩜ͳ�nՃM��[�HV1�Bz�Zm��#�+>��C��yO�˼�Ae��8��7����Hao�.X$;��e�[��5�Gk!�V+���gA���9�	d�4٥��i/�IǊ�f�S�:*uT̉}���q[������m�Q�������� 2c 	>5���7�s]����#����Zn
JV��"h�gvPN�
�"򺿗�k���
K5A}@9��u�f�װY�=vw�`�wvQm$pc�PY��a_���oYf���V�&��%�PJ������Lu6~��o3T�Ǡԥ���r�v�]L��l���j�`V6��$7��?�8�+ye��=<�
�J��x�h�~Y��$�B�Ln/b�E��Тs]���<�5\��ʶb�:�*��Cέ������W� �f�hGa2�� �=�|�T���x�S��P��َ\
�MtY`z�^�&^�D�����d/� ����!s�	ߋ�q�.�W����Xm�l��E��f�Xo<{5ܶ<�6�R�(�5��?��Gc���-p��_C�^Z�?j#����Tb�ڍ��Dd���7޾��V'���~��'���pj�9� ���s���:B��\�=�HS�Q��76zF�M���WÚ�6�L}��Q���Z�����nAi� ��07w+�^AalK�w�.���5��T�8�B�����g?����:����X|��ؗx��N�N�/-j^��COf5.��A��i�疼��3$g��]�ѫ[��O�8����(�Hg�ݣl�0��,�����"z瑞G�]�g�����nƉ�Y��C �񨍿l��4C�ը�	6�+���0ѷT�5���2�xp=��*os���u���o����X���>�1ab?q����5d�W��������9�&�v�N^J��1��.�*�*��I]܈3J�l�;��=�1� �}�F�Pxv�C�U�x�:ߠw�XV�?��y=ξ�m���&�i|�P�]����ڨ������ۼ��sl�]�'��x/F�}5D?�æ���ҪO�&L��ڵ��L>#�4J��a�'��"Ѯ�%���s���߄�-�g���x�_��.��o�a9#�T;K�K�!:�S�?<L8M��68<?���������/��]�ێ��UƩ����Xp;�����C�ި�{�t�&����8�y�H�E�Ba�Qea�K����i��g�gQY�����ִ���P��B����<A��;����\� ػpcP�
�c� ���aPMe��C�Rf���}Tl L��,A>]w��E��VX�^`��H"=�T:LJ��0k�aP,�/ б��|h��:+�\P��z4�|�,0���f%��	P�%"�٫w/w,D�5x�;q!�w�Cϐյ�|�����>2���짿����֎É�ප4��n�5O��⥫\~)�!z#U݅��GI]��D�����cT�-�NO�m�c�SXR��^��JMM���Y�����C,�ky$����g4Y�$%"�P�U��'���\�Y2��,�����p"ڟ��)�!�T);�~)?���k*⢣{ݠ���,�a�s�Gz��|�^��>���)2����:��ց�����������Tg��f;�7;pO��K��vh���EUJ�1;��H�b��~Cǯ��/�^�&�w}J�s�+mh��$d�';L,u�%yihՕ��<�	�T��<M��Sd0�¨K_`m�9��~}�ϛLD>�vu}�ږhxb8��PR��5�\�4��C 3��vk"�q��W&�h��O��ԕ�w�_RF,�0�J������W�k��h�S�S�s'�����^+�MX�����ǵF�Ln��lܴ!и3��ܣo�5njjR1�����1�jo�q]L�pO�㝨��&�Ԯn���JK���8�Z���_k]FE�(��>ܾ��$��ח�ä�%�������BTMU��0A��YI���Ok"]�����$�/7�@|��<P,���"�T�g�eeP/Qu�l�*�JW+-�<4�Gcm楓V�錫x��=�v����4�x%�[BJ��ӊ)ɣ�R �ݔr����"�������Q�j�#
��3j�+g�{����i�V��"p�¸	�V="M_'p9U�z�Z��j����@�B�Y�\v22h���Ͽmak���6!>?��ޒ:�تȰk9q�����EQ�k:�h�[Ђ$���S��;�%ϼ��4z��4L0}(< '���oC�<#z�,W���Wx��Y�;� ��.A�v����<�'=�!~~_$����L�9�~�����Ff�`Sg6��"�a�a2�p\�O/+�����	�2�{����'�=��/�6?��5�TH���z3�E?��uUf$�Z �H;��b�ƭ>�Z0��Q�
�䆅r�e����&Ƚ�.��'e������,����mA��SD�fj��XO��d|�������O0����޳��j�����r��O8)l��z 2�_�B_��Sl��=�LU�2�IS�v��qhy��,bld�lѨ��lrP??��������cj����.{fr�v�b~�K�d���d�wƫ0��C�rs;�f�B!��;-%�~�����㿫=·��nZ_^����jEJ��e�TV�
B���Rl+�1�L�G_�틠$.��yz{�^E+����0s��o��x�����2�1�:+�Tݕ�Z�}+=Ƭg5��E�8Z
�q���ҳ���,l�.�kB�-'�ř͞����_��I!�/6Q3-��Ӳ_;����fVIz�V;����Q���o9�z�5�y(�6�\x���|W`ƣE�A>�}��L�.UPI�:����UR`.B"�d:c��F��
2��*���}��(�V�(��f��+J:~_B@�*��&V�bj{�6#�yV��P $��0"ۘ�FDΰ���=�h��琛[���Zb��0
^h6����9�Ų��i㕠��P�R���g���I(i�0�V�� ��6�>j+�h�~�!�����d����|�e�pK�Rv���q�H�%��<��<��\Z�~�v/X� ��"S�1��x��!AKX !�Q�{A�QXR" ������I����c�vv�>�"+C��Y!�j��5��g��\:��AZ���k։�LsI�Lg|�.?[ba^���۽�)SM}��o�Xd����Ìjr�"z���b�@�y������; c#!RQ1�WPl��zme@���l�Λ��������;ޡP�{A�>�H�Z�� L��>;�ä�Bw��
�^4���l�?��|�Ǵ!��1GE�Y+�g����x�d��I42>���1�C��Ç����hI[�S��J/DH�V\�"k)��.m)��as"�oG�����@q4K�[���m�)[��X���)	Bt�̜E� /��s\ʄrO������d���S�=V���j�qF�X:趉�~����]�~���]�A�ڱɃI�=���P�1� /�oڛ�&n����
�)�W�qK�GY$o1U�W�4K0UZ%4�|S(��uєif�%#4+&���#@��<�͙9�����C�n������x�'��n(eTs酂�|,J��:�����&��Y�yr'��
��w1 ��L�@@��[�}$���D����V�q4B�� ^C�F'��K��q^�ܫ����[��u��e�\�V�<f���},C-%�����ū�W:��3�S����g�>��Z�4o����?e��f���K�[n*8X�X�/� :H�r`4W�+�P�{^�o��(/{WXฎ�{IB�i_,R�?6�����Ǐ�8�+p7�@=�R�&v;��J�>��~�� ��G��}>� �*]���N�%�#�a���Ɇ�v�7�)����HP|�"vx~^�����X���H�Q���^t��IIb-��}>?�l���C5M�`��qէ��&�{�*�ؔY55z�S.ouUyV�0z��Wq".1W{���{>ʏ΄u�y�^Geh����\W��ɋyi+�m�+�Ǩ�EC!�YUs>��!����!a���
i�3w�������I����ji����X'_�	�<�d�D���#׹��D�Lz�����IA��7C�s�-9\�L�^��fi�����UR;�q��F���	<��zb�I	���w���O��0���%ϰ���v�=c�^O��=�υ�j��V|@�/��Q��F���+�uA:_�c�g���R tr4`9=�,E����]�����ь�3�)^,vG��X�gV���+貔��K��ʏ�[$k����~*��<;S*^�k���?@s�"HI������V��7 *$gQ��8L�s��ĵ���l��<���?䦽"�ؗ5���u{����H����jE�s�Y�������*�s��Zl�;��RD{������1�ֱ���'�/Y�	�<?^�#yS;m ,��mOn���XlWC�z|)Ѭ�}@X���STX�+�U���}^�Е��{�"bB�݇؜Q��`�|=��Eە$M6�lO�ݖi��3�Xh��Ɔ�Ǻ���� ��fE�v�qM:Ŀ��#`];����|���U	��+��T��  �J� ���m���KB(�?�׹Z� �G]�\�p�����g$����3a�/��̃!g���Bv�׌O�|8;���;:�,�c[����j"=��� I��J��6»��|��7Vho)�����
�[�Ұ�Ӎ�O
��o)��׵�:��wAtE�a�&b� ���kD��e�fR�����Ll6 =���k}��DzC�,=�g������ ���}�#SSŎ5��̃�;g��"D�~��ғ������>)YNsfk���Ѡ�h"�bI,��{�Z�*��q�vT9~�H$3�a������Ҳ7�Ud�#��i�IP��fe�o�R��J]x�ݨNx�eM�FAQ�0h��7��k���W�"��=ۙͨ�kOM��n���j�K/���GZd���f+bc�͛�S�&@{��-�	��`fr@��]ZXȦ�¯8==��g��鈊U`��uR��N{�=�O~☂TME�������S��U�0�`�T`�k+�d8��������V��{�Շ�-�5X4�A�o���Vn

�q�FM�S+���yPd��@Juz,����o�	��X�TB[�=�1�9J,*d��(�-@����(�0o�d���EsN7��_-�r��BšGE>��$��l|������e;4�z�2�y�W�����TE$Y�xP�W��H��]ݲ��KgF�]����ۊ�rي�0���6��A|���1G������{hJ�[�`���vo�>xE��'L�g�K04��v9��l�����e�G���ŕA�5���g����5ԽT�ۻ)�DIi�Db���f�)�`�{��O�Np���R$���^��N�dR=ƥ �b�k(���M�W3z���EԊ#Ŝ�&�rN�V���3�ws�%  �#*zr4w�lgOhT�>\�ē�s/���ɢ�^P��G ikLQ�}��d.�i ��< ��*��n4�����W:��t�x��m%��.儭 � w ��bs]��+࠴��ݯ�ǂ@�BD˿�vkޠa��#���[S��뮔�BO�F_G����$�?k��0�5!&��5ࣩw�v����g��ڡ�?�ή�=�Ѕz�?p�Jκ�B-�9ˑ��N4f/j@�����dh���m�Z㢾�F�='[���U�͓�����)��//5�7�韋ҩ�zӺ|#g������G�Y
b���,�b{��^�U���p������L���H�.�1�ȅ[��p����XE�Ο�f-uqk���9����}�I�<%xgM�svK�(�hgB�]6����v6�db?>����9m��Jcl��< {.g�TQ3���"7oF�x�k+̸��v�{�	-kȗ��B��g�?-A	�M���
�y�_�w�#@e��l�OO��h�h8r~=D��x�\� fclD��(k�t�xyw���s�S�*�
d}r�:r`�{ *�846�J��R7*cF+_�,�7�N1ٮ��Q,��y�9;a'���L�@BDw]�t�q_���5��EI4T��!����B
��V
��s=�69j+�����a���a3��G2��C���ё�_p"���Xыv�Pm�4���J]C3���Q��>g�~�e���s���ܰ��Q�U�������bB��{&(.��˃�WX�K�)ۣ9'4 9B�-0�|�ǳ� �|t���J�A4�������3���٥��:��f&b�����){�+���l�*��Ymc���C�t���b��>CZ}y�?�/I?�C� ��&��� p>	�kO�=�i�b��4Q5R&�;���+3�Dks�J�ti�n�F��#yT������3`^�牛��֨)9�=���:M'/b�3��f=i��󰷺:V���s��L����Y�Ă��2U*�� 3&r�A�	��R��/(�m8�l���!��{�g�3n����v��n���Y
�=���K��@8�?��a�ֺ��[��χ͖F�������Ο�y�<UK�>@N���u�,��\���5�D�ϸ��P��;z9�-6x�3-�ė��}&�dӫ�!d����,a�ޠ	�����]�{��z�Y�M�`��y�����dn�ž�љ��#�_f������r%Mk����DʙzgZ�Ps�Q�t�J���[c��Z���m+���Gs�׳���ʃ��a���"rK��J�~W�\V��$�91gϴH`~��
�Y['��NN�n����vqr���
m���8���c���=�a�F��?\��W���x�!��ST�<���p�?^OKF�y�x��\�YG��B	<��q��^|ZI���i�U,��L��Eq�;��;��{�#�d_��!Ò�s� nɲ�@�b���QmV��l*f"G����"(��Fb������6�~EϹ�R� �L�O��h��S\�Z\����gk����=��@�ʊ�z�E��[�\�A��+:��������$��W5
=�����M����Ua3F���k���Q�A����c̆o�1`��MԮ]+f@��U?��!Cͧ�G��|y:�ją~dt��i��b�iޚw�nMI`��۬��&h��1��s/�	���t���,G=����\4{N4�e#%�C(�t/���g��f�
��1
h�$���j�6̃��O5��7�4��LSR�Z��a]v^^ELT��<�k(4�X9��kZ,��_�[���_b2$l:^f/�=��IIyr�\Z�c��*��V귭��v�/֪`�/C�kK�����q���M;��An��h����sf�$e�նI��W��Dx��?��f�K*]R<��A���޹k�Vm����YU��}B&�ڕ!<��L��9�O�S�}����X��ʣX<�J�T*T2�`��/W$G�S�[Φ;���3U�J2���B�k��k������T_OX�rMU%���% n*9��Bg����3�M�p�HF��)�6)��^���>�,٠�;���2���U����� ��JN�{�"rs��U?���Rg��g�n�\O�Eث��7֟n91f��[bX"`&�c0���^۰}�\q�:s������-+]��e�"r�9��&%T����v�o�
a�+�G���j5[�;e�A_�æݡ��e�zۜ��������S�%*�����<�(�Q�4���i?c|)Bp󧉉��4���~�N�-��y �0����S���;�[��<�sr*	����3��k�F�X͕������*�X��T>_��j�;����fN!�a���GfPR��^^��^�~\��{�kRr�+�J��,�t�ǰyNԊ��=37L�估� W�dpY̋�]���ł�Z��;�cV߷��ci�nE�)��
c����x�>%A�$c�S��b"n�j ���M'����������j�����u��"�J��u�@��C�����b�z�s_��W��#���vu(�f�'�e&�\B�[�ɘ�������{V�������LC�d_�C����5X<�YM�lD:��v�8sFb[���B��Q��xr����T_�s&���n�S^ޯ6�-��4���&�=#K9���$O��%�;��v]Į����ɟ��g�s��Ν�GJ"�}�3���{ɀ�yW��屿8�l�?-�)T�L���܉ wn&5����7�]kd�P�}����r4�I5�<��?瓶�<�{���M�5�C7�3!�E��+��R�aE�����%�Q�%�\�1x
H4��w�쁭_�ڭx�u��J�?T���*����꛼�U������%�5j҂�&�L���L ��)X�;|�
:a��*y�Q����p;���_�a��7���(�ϸ�י�d<C
��<���qGT�J3���`��#�æ�7k���o\o�]�oշHs�&#^�D�O/=M�|���U�*m'gƌ�����w#H�5��^��gʾ��6�ʋ�^�>5���z�v\����Y��@G�Y	I\��N0K��`�����T�I��������z���f����@u��ޑ��"](�{)��[����٫_�Ah����Ŵ�2�$A6m�2F�R��ܭ#L&���usWo�O=cFT�kUߩ���^�A��9�*�������z9�U��!��(���7/9���|NU�1������><�(�S�:N��RgW�i�����Y÷���)�aI�����@c���ـ���syx�	���Rm��D�d��/@);�z�U�pv�$8j�/_���[\�11#�x�A�axga��l�z�1ccE�H�h0�����K�=b�f��@ݘ���MJ�GV����% "&���,/fZĪ=/�g�����Kt�O1�]��9��U1$�r�m8�F2@�_������\���ۇbǄ��)�c��?��x ����-Uc��I٤G�X`�H���ckt��o/�Q/,����^]��L�w,NK�Z9�\1� �;�Ub\�?���]�/�Xyj
�8���8-u	d)����~V�&�wG�#�D�<]�G�öt�i�۵I����mj���<y)����'ܮ9��^��o�	�����ʖ�򟯢H�Z��)c��G�Rrե-j�W����9e��s�K�P?@L�G�X��E35��C�]��+X�%:�����8�����L尩X�u��i���ˠ��m�e����^�����k;ӿ�3�I��&����5��=Ch�V��6;��6o�6Y@^�nT��6���-��[z��]����-�']���*y��I6b��1�e+HV�ԭ��&:|iBDσ����z+G�`��	�������M#�׉e�'J_���#5��ܬ��?U�j>��k�#�Z����ʍ���re+ѹO1%K,=�����+����N�]�ȷ�[نު�xo2��]?mB͂u��t���.�»L�0-7��N�dJ��"F�0�B��&k���fIB�縲����Dw�Ȥ�/jq��y8�%�\��a�Lm�o�x����-��(�nn�K\Z�����Ȝ�	�v�G݉9�PC�<Q�aⰢ�@t5+=MzP�,N7�M����r�pP6W�"��X���_L�r�k�Z�!׆���H{))W��3y��LF&NҠ�<�.�4�^�|�בm�3��*O��hF���B��a"��'���(F��mW��w�~3U��,#�ǛXxk5w����ǁ"��]Z�"������KQ��W��A!�!���^���^����(N���}g�f��U~K)$l����A�w�m����s���ڕG�{���Ʉv����{�Bj�ƻ;�>����a�+x�5��<��o�?�v�@��l_��ƁJ����P#��CI`sl�[zft��ď��e�$��<w����__u��D����f�	�R���&cI'Z��Y�ZV����ż��~\s�x�߹}>E�Cjw#:e�i��8�Qj2�?E�K�n��᭜k��ϊ������O��7R�wo�_'e�Ժ���}:��5,@ޔZ��i�a��,�~Tg�FJ��b��&�hޭx�qE��k-�%�]h�G�RT��y��B|�!�o,��p�B�k�M Z��@s����_k#u7#0>)�^r��
n�{T���R(�K��;������EY�9:��殆���S�*{m���X~k����b ����f�����*����KJJ�L����x˭�J�'8`�ߛ�A:u��.�����s8��J��~Z�s34f�K���eJ��RY����ӎ�sGy	PˣU%��enG���6���c~z�b�J���g;%��&�φJ��<����V��P��y)�f��?�x���s�	-h����JW�מo�E���'����ѿv	A�媌OQ�;�����jI�1-����p�+�f��-�^vYy:,�:e�#ŻP�.����A�)��^���Tc�w���]X��y%�n��ܘX�\^�i�|޷RP�P��n��`�;��:�u`��w�.�@�D��`������v��Qa)ysU&s:-�O��E�Q�j����	Ґ�>�9�@��0B;����*��Y�x�,'�y���n~P��Kͱ˷/Jު���H��^�=�(�g��4��<M14��;H���@�h�R�~�J�b�_��"�zn����+�8�D���M�}��O���m*�@"(����Q�;kJGT���C�4���4�&!]�	=����-5^�q���5t����jF��a-i4U���	˗�o���cКLc�L}7�ŋ+�w��p�^�'�!N/zӰ����D�TQ���!���;����t�(L���ň�%�n^E���ն��vb|R&�6٥a(�E����y8vn��k�*c�j%ѕn˻�,�גWG|ٯ��U��Cq4xZ��BC��a?YE�mi��~��p��]�kep􁿢A��1u�r��<{_���Ú�<�73�=c���l����-���qE	wN�N�sh�8��Z+�(�Q�}�*>�^�̣���{22���a[Y��kQ�,.f���A�"��:*����le�<���V�d(�׵�sZ�z��1�l��9�rb(��m���c��v�@0��A������옍�<v"R7���zbX�3Ğ�)~}X#@��0�jV���hz��l�k��`6s����@<�!�nZ��N/	�������\j�t�z�F��n̄H޻e*;y��r�*��Fjq^k��C�%Y��e3 ��*NV��;��i�em�j�W��vHV��a�i��i���� �!�h�-թ���?(���w)m�7 =���CBӨ��	C(����W˒�Q����}E.Ve a�Z�����*��Uai`"�I"�$@k2]��V�e�L@���'�R	"���4	�:����]\~�Xm#�h'�GD{Y21���*6c+x��v��L�80�UQp!�"���ǹbg-�1xB���L]H���-a�P�䙪;sI��cƍ!��0KA�-2�:n)��ʵPa��ؼ����w�]�o�8�p0���)��;t�GH�7q��+qQm��Y=���|���K���hC�������a�����л�ب��7�3�p�HĈ�e�Waq�-�nW�;�hu�k�<��1����0,�������=�ݧ���4ڶ�I�ʓd�����F�&�g�� A�]K
��w<�ͶX�08%�݉N�ʻ ald(���$3�cRݺ���"�z?#z�4#c��[%|ޯ�F���Ƌ�<����S|�M�J	S�r�6�	�Z�/Jt�E�o����47�� X��M��sX󁹐��	�B#����I眀�g�X]$��5dRb��Zn�t$}�N���C�Ljs�tr�Z�����w�:p"���Y�3X�>T 6���f���ROȗ��]�H���vU�nK�w�M����qBZ�?|�NÔe3oЗ�
��x`Tݼ璗7�%O�iхr96F��N���s��q���OJ�u�s8����ޮ�9[����r%��>�߽֞{��;�qRT"e�:��L��[�P�I`���d�"�����,���-{!��p��TYR��Z���2'a��0`��ӹL��te>��}3|��^� �4k�y84#�BI�Ϛ�&����X7L�̐��9�5;���>6�1뎢J�] ��5����T�� _�q��.�v���Bߺ}�'����Ng�\%o�u����X T|�����,����S��3BW_1��.վ������Hf�����F��.�8�(����R�k/��8��_BEȘH$no���ʾ�6����ʰ���m@���G�;�C)�)AJ�;��!�C��v�n$�k�;���^���8^r��묽��^�Ƿ{�3��Z_��ûhˋx[P���;�
I�Fa[4�/ۃ:�`��n�84F�B�ڵ��x�����V!rž���Ke' ��Z)���%"z���k�֑��u�������͇G&F�^�Zi��+�A�_���焜F�)�(�]�v~��Y����哊`b|Y�������vW�>���T� �)�O���W{��Ŋ�ε;����GeWヂO6���h��?��O_g�&$����*�c����w��K�Ƙ�<�8'�>e'��Ԫ1̦-��2ٱ�%v���g�)<|%#Fr�ۥ$V�#���[��~ڑaJo��>�g�Ye�٦�q�W�d	�~�|���|S�č+7 K`�n7�
C݄��O}^J����A|{[ڛ�ޯ�H�*��;r�b���fGU�<��2�y�C����o�f�a[.��ݣ�Zc�}N����`:�jsLv�jE���褷��3J��:��wM���L��D�p�]�9��ͪ��q�^�����Чmb�#�T6
��2"���&�R�� ����U���rD���e�-��Mol����oG�Fj�|'{�ߢ@�7p��Ch*C��h�r5��f�K1�O)r�L!Č��K��		�L�2��8�ؼ>G+��L�+�F����x�����O`D� ��D�6�-JR�h��=+T}��#NL��/��|Ig��Q�"�XH��GsdL���
9+C �X�i�R���,�mx�K2�NP�k"R�`���r�·����j��g;������
�RRRmw���DW�D!��RU�-������t���W7R�X������,�����l��7o��ĂU��u����\ O/+��n��
iR���ڝ����r��8��h���g����`:�쥏�̠6���"]�X�ו�(C���?�;\���8z/�f�X������ub���i�k ���~���l�����8��p�h$�RTûI��?����o~������������]m�@ۗ������I�\�a�\�\_�%W���NWi^w���3V�̟K��ׁy�*��M���#!��u�u"����;ۄ�:�����B�S��S���W��g����H��E�Ҿ��d�pb(����MMQ�Y���k��V�ƿ�ao�do_ޡ�q���ޣ��k;���s2X���h�k%�|�C����J&a�x�P��>�f�x�p*�����Zk���4,N�&�k�pg\�,��V�Щ)�?:�f�x����tc5USV;��t~	�~�S*�X
�j�ڦ������ęIi��	���/��]+Nt�0t�P��r��+s8}rW��G�6^Y᚝��2��[C��O<0�Nh��2D���:�;���9ܸD���*3
%�KU�[WW\��)gn+(�)?ᇔ_U�(�2�J=�K��Q$n$��3}q��G�F���{'���K�����T���~,[`��C8������fdTT��������
/�U�$�	R�=Ec$z��T�b�mն�Q�&�̮&uc���t���� 2%7� �����W���脏įY SL!����������t!JQc�~��E����"��<@5�$U(��w��ڇ[{O�����!�و
c&����=`5��K|�� `O<zxl�p��GK�w�_c��-�C�4?\8�����S[����h�� �C��)K��k>0{I��|'�!�;����@�\8��@� '�?R�#�d�n�
���/*0!~��[��ÃcȈQ������iX��DG�:`b���������� IG
����0�~�h9�������?�ATJP��o�HF� $����J�����g�W�j�'D��� ]��o�+݃�e�#�*��\t�L�* h�����GE9kq�߿����������'��B,���?���o՘�k�|X2���%K�FT�.�������R��Br3�QG��Z��X�k>DvB,&��.��Q/����j�A,CS���q�Axp��7�1���aFħ6�ߍ�J[���7��Ӷ��w{���f��u�+U	��G�T��������� �n	�h���m$_-�&1�Ě�1>͚��cd�2�j�k��uY�'I��{5�w�=$Ց��,)(��

�U7J�\- �02��#$9E�:�vW�O�!���d�A`�h�:�Z���ħy�R���^�k{� ��޾��2�e?|� ��ٹ<�gaHк(�D�ց��"/���b8�0 P-�����aw�ſ:::N��:N,��ߴ�X���<�!_���`Uw���k�`sB���k������[l6X�Λ�	>X�7�%%���/�W˜י <f����P��|x��U� C�БckH:������6wM~K�� })Z����Q^�M����M^��h��We��&�T/n��G%�"i�Qe�)nsrtտxj@v)�vq�7>�&m�*��jCL��������}{���}����:�ɪ!6u%����x����CwZ�ic�W_�|_����h�%����Y·��(����>�{�4|.vp+8>'cd�r{���Y����u'Q���[u�>�ܓZ2S����2�Q�. H~�˂H��r�>>��ap?���pLD��+��������՞"���0��Yh����+?1	_Tڀ�hSZ?嗹~L&XM��)���\�������)��Os4f�q�mB�O�G'�����+&!?��/�iٷ� ���<���H��:0��>~��_e����Hk��񊧌�e���(�V2~=gUR��N�V-���e]�~̹��W�+��M7L��:f�b1ʣ'��ГD��W����:���/���JS�)�/��
�H�I�/�y,��b������>���;���V���0\��؝Ќ�T��}��L#?�.@L����Y��� o�LPz�idP��zX���ib�a����'Ϸ��MYoE���q��76�f�<��d���9�G;ŀ�+�.T���r�w�1�G�H��CȠ��tᗹNh���2�{|��r�.��1�V~gS�������v�I�H2��e�Q�tp�ꠁ{�{�b��"�����tI�!'JK�`�	�K�Q\���;��2����Bl�nZ8o�̒m���0MX�����9G��&C��֖��|�8V e��3�Ymtm�Z��{ӣ��t�V�M� ��?c㐑{�����P�!?ϡVm�����(���Q8�T�3k�K ��T������|Z��i�Ǳ2���:0�͑�����L������G	�DO�36'?�� e�u/u
��兦Sc�+�͟
�1��Շ%GE�*��+05.��� ���Eh�Jyb�{���uAd<y�_�z!:N"6����g��Ǖn�U��9�T"O1Ee����q'��g�68��>�x�6�_����h4��<s��=���7��kݳ�G�G�uG�	��;<%cmo�g�<��O"ֶ��������/�m�5= �P�P>�K[��,����X�G�y�5:�`���r=�97�Cm6��S��T��}Y����g��k)(+Fo��R)8l�%�%����3bRD��%�%u˔vyz���+�F��r> "2"�"�Td�:�Z12���7���nT����r�V��ԏ,��l),�I���tq �T'��v�'��\�����1W:R<}�<�A�CL{1E-ʤ�X�w��lᝑ6;"H9�x�b�Ա�w�7QU�	3�� �Y��NĿNib�jԫ��nU�#$�%D�i �M�����݌�;��"�T���-�EW?�Ўkb?�y%�?��ÀK��b���o1	<�5)C�H��o�8���?Iϕ�7��
R~
��z9��I\�;`�#a�"�`�_n$�S���:6u���,� ��]M+���A8��/��:dp�����-��ħ�S�5����p��3��Z[�as���_�jg�|5�#�K�Qp��;)�Z;�V�Tc1FREYA���MbP8`b��w��nE#�\_C��v�]�\ە����>��PG�	�1~B?#�K�9�Y����~~�L
bc�X�e\qi9B�uʍ���}�8Q���dl��B �j��f(�ҍ"#
��ճ!ω՜p��w�.��~�a	}$͞Җ�#|�0aV����Gg���\�7b�T�0���4�?C<���+�E�ҋ�i�VٽYZ �ur&xf����|�l9d,5�F"E�CZ��\��C����f?:5�m��mP��=����b��Iq^]��T�kFғ�JU��n�(:��mE�x"n�\����h%��X���+��v�.?��>)�VH���o4��o�L�Z&D����|u����J?Vk���d]p�'�rn�T����U!��Ke�M�Ǫ���SU�v+��%�np�{ȫU$H\|0FA9� 2��q�3��B�
}�O���Kf���h�00�ٷ�����\�0��?�V��{��>����\ҙ�hʮ�06y�$`y<�d�3���}��;��3������@�<4�`�$��xG���t ��:[�_?A�)*a��bǊ��E�fI���HxӒ�ĝjJ��L�]i���I��pfo���>��.��$bӡ�rG��/}ml(��*���@ne��1�M��7���\w�T�E�=܉ !�����K� ��-��d��8t/5 Pt�+�c��)@���u���.�%W�]
���x��W��$�2 �]8mb*��-|i�c��`K(��'A����j|�P���S���g����+tj��O �&Ig�c�(Ň��7�r�fd���Ľ0�y
��{�$#�����Ⱔ�X�ZψS{o�����������ث=*駐��$���V�/U�� V��^k����QA�r�T����W�h(H���_F���w����H$9�䏯t�R3�~������O^5����������Q��7�����p�b	v����� �%��~8+�w�>4��|�� H���m�u�� ��6x,�ܳ����_��|�@%�e^�#���^N���8�DJ��˲�U��E�r�� �o=��D)�"Bw]e�N���:np.DRH�3b2�EɚZ:�c�?�~��`�J̸�5�E��&X4�83;���l�M�2�~��Q4͖ؔ���/�^���D�L���ϻ��㸷�9G�-2<���B��Bb�_�>�s�Ң�w�E��	�u���>�&<��4�'Q�˴Z�����'��	�Fb��Si6��t�6I��^K�" �3)#�e��I��i��JV�Q�����,������.!��a[�����#=�����x{rhP�_�Cyf�>�XۆniOrC�ȱ�v�Q_
�~ �_������:�-	2� ��I1���	�>l�P=���Y�v��n�t��"�a�ܾ%��υ��̂��ց����4�ЙvJ���Jhͱ�0j֐���=����u��ݴn�c)��[�Eu����X}�z.���ط:0��c�C�/O�*K�����VX�'�=J!�0W
P8�jV)n��6���q�vj���K�>ˏo���73V����GSV�Du/.v��TY�����o��i$lX�K���uJ[a37(CԺ�m��~�[e�!0���c܅Z=�|�Ǯ��:�`�Cj_��� 	[֮	X�q*s����C�r�Bm�O�m	D����tnas��KUG��@�WGƐ��"��#C$r `vJ��sG|��%	���>����6b�<�o ��mpD2I����X}"�8��G�gFk�Y���=���1�?�fz���0��=��p�0'R�N��� M�`:��=_�c��MZ����I*��-)��@�Qwo�s���;����{�5�>�Hm��4�;:���ƒ<s�@L#��M�h�#���5V5����/%Ĵ�/٫oZ��l[��H�4f���/�W)����/�.�����(�r�:����iA�^�t�v������Mk�^���ǃ$�k�$�CI�7*ui�v#��qOQ�4#ӝ��!չē3"<��8KN���  z�>��k=��'V��I>_�Z���bʜi=M�I➫�[�"v��y����2���	�F)U]��@=������to��!��%�dSxk��r��Uq���Hfzi�\vC�O �[MY�k�f5��K:�p�l���#��J��������r�Ȓif��i�gb�p��CT��+N��S��p/!���]|\R��K�����[�|��ҝ6��)������wc��Fk�3��Of����U�^��I�2Tf�W�^,rX�no ��\0�#I�;��E[�p�󖫩u��{�����r�qH��:��(�3���6�t��t��i�/Ru� h~򳁕�Ĵu������m�4;�iG.
��"�'���k��E��®%Z
��=���T����u;ZwO�H>c�HRw��kV���)��d��38ͷ�zs����<�JP)D9�=��!;��n����<#]��e�|t����@r$��x:�7G-��d�,�!��۶:�ݭ���5�V+	���n?�#��<�(�L�d�X�{u��.?>�;;�>)#�)�X�QW���>8F���K>:qg�����?�a�羫v���ka_�m�s���CQ�����c��ٌx �R�,�x�v�k*�>�z�K<�%�������D5�� ���~_d�� _��M����bZ�3��1}S���e�ǿ9����:��Tq<�aP������>�!�$�ͥ��z���T��%��D���E�X�&BRآA I����b3�7�U�����D�� ��?��)ވgޚ�%�΅v����p���|�MA�t:��׊���͆�N�M���"Nk��b3/�㟋�����ƍ����4�\��r5Щ���\����fgS����%d7V�V/XW]w8��7�tu��r18�n�my�N�qU�#��S{#�Rm V�KiB�²�rR��~]��&;��@��uX��r"J�J�5]�D	�'���a�s&,r���=B��*�;k�������-n�z.�鬋�2W$�W���rr�f$h�p�����'R=[&)Rʓ�ǇY��I�?�*hl:Y�T{�ѻԮ3#��Cgt�̶ԼQ^,�i��ٓa��7r���<�J���!Sx7��I�o(�N8F��Y�>�5��~�XEh����_��a#	l����lu3� ���6���h���z(�XB}�է^
j7���<w�͏����&��@z�����y�,4zn�s�4]�_�.LJ���.y~*pjc;4N����j�����f���%�,�(B�.��|7�\�Q���2Gfq��deo�r02��������6<��n�E}��`[?��0c�8Ϳ��QeFJr�)�r{�iyP���M�����ak8�����]���Ku�F�񖞂�~�]���nsF~����FҼ;�+6��OP�tc8�̘jcg;�VS���*V����d�0�Ob`J�Ŷ�v%�.]���S�K�"�qAsȤ��i+_��/��;��H�?Fw]��1"爹�D�f��������iqt��"��«#�!\����<�%��`TOC�ѿoY�O%`��^B ʑs�1Q�r��l���㎮� ���8���~���A��[�), >�3�V	�,D	m%=�o���}��N��\�J`�w��s�a��uIɘB�l>��IV_�3/q��K����+�Xn������#)�J�9��M�5����= �m��n�S�={Qێ_C��X�������Bhs�}�m���Tq�x�iryTv;2f�w?#CBos��""DP~e\]I/�o8-ߘ~q��my��92E��E�񵦍'����>8"xK��:N��-���&ֻr���}������U� &D����!�R���!рpdD�I��E ݢ�yؔ��岡��Jb��sO�1�<���~T�E��7ˡ��`a-\;��x��e^����N�y��zd�$�4E�2��ޗo�CM�o[�^4�tf�g�gѬIo�p��y/�S�����Q{J�R�Qǝ�Ǩ�d_����6�����XF��ъ粕�_ruv�
D�n���cj ��g='��G�x~p���A��w^�T�U��(vg�l��8̡�cf1�>|h����D�h D'���s���"O��~��/N�m:9� Aw>�(�q �	 ����6I������Cǒ��w+���Ѱ����6YHZ���1����K!���׿ˠ��Tr�����P�IEH�q�q<�ڠ�Ы��kM�W�o��kh�o-�A¶9_|t_��Z	��2{;W�Ap�:����[�_�4W�������^�q�+U��{{����q?&�۶Z5��3�Lk��[�c�+s5��$�2)q�{��6��;���˄%��a[�� T���$���>��0?�5���O4�j|*|�}f�D,w�� ��ִp	����
'@G�C����:�h71I�� 6ع�L<?nS���LM�OM�K\��6���^�]h�,8�%.[��Y?����R��	y�����W ��;�r�	��x\�rÌO!���G���{ �/��V�cRF+�&�T�&����}_I,i���������b��Ίz׵%�>C����t�4;�N�ht��jw��ʾZ��ͻ���������?���S@t�s�\�}Tw��:]8�{ S���/��8��H���zy'���|���u%������ZQ/�#�X������g�ctӄ�&0�����ʉA���ZZ��4����n��d�5����kQ޵G�]�]�z�RQї�B���(f�G�}����Iр���T��n���Kcw7m?��f+l�	$nf|��u��1�ea�y�A��� _$J��!g����=���,;gq1_K�w6�{��y��ִ3ֹ�c��+�QtA���N;K���}�����{��yߏ,q�b	��d�^6A]��K�8|�f	X��,�̝�S���YDK�|�h�,�w�)���	5L��3#���gQL�|x���	ؗM�d�d �
/�}i�v�{��x����}�w\F-<��3 �x഑&�h�	À�a0��p��w�BS��l��{���������>��;Ã���Uo���Z�_��?��pW�A���p��,^y+L�9��i�r��IU�ސf�%|.:,@��X�`��[�MRnC9�����£��-7�\��B�/ޯۘʛ�$�%>�����+�-?����_l��Uz;�R�ٽ ��^��yH����7�B?�4(F۶���^fE�{Ky���~����-7�B]N/�v}W����&E����*��ŧ�Sz����iW>���`�Km��V��I���o�A1��4�[昻���Z�!i8M^� <����E^!}���%���6��W��|&�M��S����?f~�Y~���#V��	�Mw	���R��c�w�s~_a�����r���Ql�.C���eK�w�h���]`�*�� �/�����h�ݶ���E�rQ�w�""��x��g�M5W �*٦UZy���~�Ϳ740i՜���t^}�bu�µ_L*u���>����sU�����)�Pc\�d�N%یK�/�k����5���>x*\�1
�!�� B�{ta)��}v,ty9l�R~G&'�0fw@��0{i��C���,���n0�T���_o?q��x��ڵ$���)$�O+�^*<P'C��D2���w6�"�͡p��۫�R��ؑ7���!����O��!*�>5��q�Х�|�¸6Y!"�d�g6�<�p�����Q^K�L-�Q�ҹk�x39��c�Z�e{�.�/�%V�׃2ҝܣ�P�ݚk�
�IV^��m+(x��Pf�=�X����a7��͵�Â����ݷ��a�F�������Z�A��H����m�����Uy����2�2�6j����!����9R�'Bz��#���أ/18`}�����2��31��9���8�?��w*���}���9	8�}�=Q�Q��ע���c��j[�k���(��G���
[�Y)r̴�0>K������26S�E��bX�
m]Xz��՞�(Fo�6'��,�AQ��z���$����f��dk�R�>����<��������G�j:8)n4��������f��=h$��DT [�S�g��"<g~Jg}��7��1Cب�����l\��}�R�غ
*e��.�/"��1W|��x��0�l:{�Zo�?v�\P��${�m�LMQ�W��z�|�3@��bs��I������AX�[���V��ȻЄ����/��wQ���i	°H���/3�x/ŗ�WK�϶�M^yK���b�cS�w�B���}xv�y�5v�/��`��s�����X���d���/�^�X�W�d��\��87���7�s�d�J�|M�	�h��>�Y�o ��S�V��`����;����H��H������ˣqgG�pF�����������M%ݥ� X��Z︩���V7��E�_����E��$��K�k��7�"[��T=�|��&&;���1N]� �(��6:��D���{@q�	K_qmSڇb����(rĩ=�h<�qr,n�+>8���^�/L�n��R��r��7��+��*�E��b'��̽=L�=��l��i$ԱLp�,DA��W���'��ɴ��z���3_5ʝ�}k���@�TT�_�� ���� )��;�}W��� �0}�{^�΁�&70���-;]�b��T���~S8ފ)0c��+-Ŋ�g
�?�N�Ά��*Yabң��S�Zƥ{����U�*|c���d_|.����8Jy��D<�@�I�U�[D����ZOq'��m�����,nz���2��|�Ǔi����6񾭏o:�����d�G�턦h9L��0���0B	���Zp��塠�?�%�x����.�T��� ���i�2M%��z�j7�?~�0h��2��w��<eQP`��aͿѳ��:_/�ҝԂ�~E���k��1�@�� �f��m��1?���O�}G�}���dQ�4i�����Mz�3�B����"�?��%�"���9�d�۩��<���@A+.򌳭�����p#�¹���\Y��+G듷�1����l�c�����Yu|6�͏/Չ�( �D~j�Z~�wQ�6x�?K��~t�rS����,�-y���͂A�RNq"�N���t[F�>��GO -�$�m�yY�&�b�/����qӎ�u��\؛��[8���7��#芶QSF"߆�>��j�9���UQ�3�۱B0�u��oǷ�t�"
y�%�[��#�o��k�>�O��`�sW��|�h���;�e�~ ����ˡuPF��3���ܧ�@�n{��v5��N��`�$@Ő�[j-�a�ֳ��o������U!	�g��ꆍl�U���s�p��;'W��d�ڝ>�{^����
�9SKԿ(!8,�����O �L��PT��߹e�P���q?�Uü�r_B�63����s%�Ν�rs�|~l�X��"�ڼ�qM!֩R!.�씶�s�"5�! �V�a�����.��j�M\����Ƒ`:d��:�i�w3XRd��BCf��O�[꘭/�żMe���r�q-?�(H�����h��8N##����(@�&��xYyK�pr7J�{�Q��1��.�Y�1�A�p��ae��z/�9ɳ�w��w�ś�U:M���>�,�|����H�.��5��|v��enX������h����U磪�K�GR@g���"p�g�6��]i9eO���_��+�W.
�w��=2��1[*�}a�VIf\�U`}h�#z,a[�J	����`x�ɑ�C�"+�Ů%Eκ�s��ڍ�~
�'MY�ID�+!wKVC"�$^�����hv6�F�Ð3o�rWr]7�tH4�Q�Y2� cg�[j���~�Wlc�݇��x)���,Ba�Ѫ\��J�^b��6���F����ң��`U�S��/3���|tt�f@�W������V�,"?�TFe�vQ��t�a�����[*x��k6����9�so�#�:v����c۱;�}��e	���%��B�hp�����RP�:;��פI"Sb��~x�H+�9��ߖ�J��t_\n�� Ǆ�0�$�5�,�Ap<Ք%֜��;u�<�p�F�ߜ�n�=�L����\K��M��2��̹l1@�iͥ	�^#Mǔ��a�h�u�����j�M���#e�k�i =>]��r�B���L�T�N�cR����%/�������u��4��W��b�,���_{2,��������{ (#�\�MGS�����%�Lw#�c�ܹm�TI���Tw�m̵��og��1�QAK=G�+�uT����HH)���bv#pA��'їC#�ܓ�8R�w�\Fy�00�w>,*��)�0�jaJT�E��oB�o��Bl��r�LV$�H/X���/�R��I�}�����5bI>Y!�>��;��6Ρ�u�j�s��ܔ�.)�jo.ο?�Ѭ/��['��H���(&��)A� $���e�Ȯ�%q�C����;���ت����j�T(�ڔ����λ�����g��w�bn�g�F�BÖ_�����q_����e�Q�7�������%�l�o/���F������U[�23$X��{����$1s�x��h����}7�gٺN���8B$^+����!]��E����?1u�4����m�.@W�,X	_�V���r�V���e��Z.Lۇ
|�����e'<��]�j+^(Yt��O-C(���j%�ލA��-���'��#��͒P���_2�C}��:|�~�j����ϵaLvQ*��l� �?�����H�&������݇�plu��E�QU�����	e���`fBt1g/�VEa9�AL��L��BF�/Ԏ������]��:�����{���+&�+<���on���/i��E�V������ٿ�*) ��R��/g����$��ߪv������!�Q��
�jz8���0"+c�v����ώ(G��5i���0��C�F�*@��7+a[�7u~n��|���}xyJ��
��࿬�}"�e�ɽ�U����!�(y��gK��ӎ�\h��K�S�G�{Eʝ�B
��k5k�2׿���+�S��P�1��@����v�J�MzE��<9�%�\�������.�n·j�?�J���U\�+�*�J�j�g8`�|�����2ں��ET��h�w�)}��H���U-�����Gw��c�L��mF�Ѩ(s�G�<���Gh�������/���E���ߨ%��2],?��o�vy�����|sQ��&k��Y`�D�4E�̐������n�����ɷo\����/�&Ͽ}��51ii�'�ә���I�8) {�=���|��ʇ�[CC�&nn�A1o9���-��H=��XM�FS^�F�2��b��F���CB��ĠU��Ҙ�$�Ɉо@��	�#���v�z���z����O�aQ���4f��K��Qi��y���'<!��l�[�r��8ha�>�t����8��������땗��E�� e~j+�{]��v���q�,�#fE��͔���$�~%>[*���T	�[�&���}T`���ׄ����w��돾����6������5.^����h�~�o�w�R	��.����n�G #&�(wE��j��h �ὣ�\��˺lYr�uxK(����oW_��۞��؅'꟨��ϼ�S>ͮP�C"���[��b4[͙�z$\���������HK<>��0,���ݩ���y�/��ۚiEC.e�����Z�v���@-}y�w˗"�AW ▆ I�E0����vd��X���cBxq?5���u>3�r=,�wu�HE$ul��hH`4��S�է7��W�_��f�mZ8XU�n���a��j�7A���șrX�	F�̩T��9�o�HO�G���T4���R�ˣta�b�ٞtq����K�)��:	@y�.�o�]�U�!l���R:���u���ŠI'm���N��?�*ޭ=�ήm���
"�*{\Y��ҧ.��{��NւQ\�[u��:S;��]���E#�Ӝ�j[`�6n�K>Ǣt����H�i ����cX�I�tY'c�����]$���`�	�큲�U�F�p��L���Sb���Cf��D�:�Ѝ��[�U44Ş���ty9'�	���ph��@8����}�'�Uy5?���t�<�
�5�����K���,�!�'z�6n��C9�fx��Z<�j��5`�1�Z5��~�V�e<�D����y��"�oYq�"��G����SUj�M�[��ށ�M��v}�����@�cM-:����
q�d[��>Xr��&�����g������n쵞��i�m�a��t��8���D�k���H�I[F�!se��<���S>r��(�@;�_�>*��W"�����uMDQ3��?}�p$���D�S�j�6f�t���E}W�U
��NK��Cx�b��*]�5E��d�Z;W1�w#��Ou=�:_���v�E�������ŧ_>�j �AQ���>&k�%��w�UZ����<?��&.�-�8ڰо����������p9D_�CX!F���E�W���'v�٘��92@(���x���%ݔ�s��ifj�!�^�9϶�ʼ�EL��ĥX�	��'�̉���*�#�6�,�k�l��Uΐ��e0��SD'�%��b��z�^��R5�e��m႐9�ϳ�*��p����:ǀ�ޝ�|;;���{�o8fۭ�;�+����bI'm�l�����TG���:ۖ���'�`3�/Jm�#Z�����g*�(/�\@Ѽ�A��qw-Ax����NQ;���{�	˕���X��#�/_���� E��-�z\��W�Ur��ڦ�v�U��O���� ў�9_Ts�q/=77����\;��Aʯ~�RP%Z�k(V_�I� -�i�����$o�o=k��J���6}�d��)v���.���h/�A�5\Q�w�I�L���?�gtx+�ʵ���?|D=��1�k^FU�8�0�ev���1r�4�{�`OF7�K�V� ��.&螸�C':G��O��>���e�^u�k}p*c���@Z�\�؛f���|�@��uJ "��<0�(΢xO�2�!(���^j��ݨ���=YB����{~S�z�
�x�	EI�Ĕ-����yؿ~w�5̌"���0@
G�F�q}-1b�X8*ۦܧ��l��¥"��r�p3�x-m����-xa���]1��Q��5�9+�m޳�՚�����_��l�j3�Ͽ��t��`���7@����κzq���S=l�q݅Y?�M�.�:~���b��tB�8�N����ʏfO3�sH�}��8����f}*�q�ѕ&�a�wmWv�gK%e��zq��\����cv�t�n������"ϨaT	4���hSŻ0��gŷ�[�����h�&�	A��UAс8��M�E�I#F�l���B��\����q�>���E���@�r�[����L@19pȦr�R�H~��G�ݻ�~��#ތo�u��-���Aҝ��g��Ļ�i���n����ڴl?�����_.�ƶEO`945٫�q=��F`���'��t�ǌU?��=zߖ�^kߣ[�GG܈�^~y>`h��#qw3È���#C�,���^�P''[ȸ>vef��mtH��`��|����J�/Nd����M9Gq��'m����d����h��8~��([��F�6 P���� y�Ej���Q�.{�����j�.}��&7$;(���4��']����X�n1�|��f��~x <Ʀ��OC b�/�Y��v���9��vA2;�k���%��*,������C`��A��_N�'�!e�H�����Ǹ���	)}�6:Ջ�m�Y���)ؒM��aDc��D�''��pGf�O�ަ�t�W�G�[ ���$L�#s�Q�e���q�����/dB�&�G/�JZ�j��CI�8�Rc�Oq u�V�|�q���tJMSH5�[X������-VE���Ry@����[�s2���v���Z(�$��{�:�ߣ9�\�*κJN=7 "�y���E�vL��ʫ,��Do��X9ìk15C��7��t~����HS��W	��h�6M:�� Ξ�WMw�����s)~g�fɥ��c��O�x1�Q�,��X5al��Q�\��n��� T&��6�N
5�����2^�ۚ�zؒ�Zuޏ��j�0�~Zۗ͐!��AN�H� Ev����%ɞU�l֦�g��������0�Ev#��>�>G𭀈���ibbb�MMq�̃&�gD���Qƈt�KV	���@�'U�}�s�V��Ѕ��m[�s��(��4ޣڀv׼%���'�SJ�%~8�z�۹T+S�������6��!#����ml�tҎ��ᑡ�,K���~��:��!�E'@���d������`�0kgא���
eN�o�;-����ב��*��Q}�w��y��9&��g�򟾅�ɠ�!�m���r�Fݣ1�ge&�S�ߊ��4����J.%s�ձ�c���[���[?�c�m5mt�o�*��_[��*���0����=����V致�e�+x�|���w�9_L�??�btpEIl�J i9��!K��2x ����/_#�&.$�	��f#��q#�fJ�<�m2q4*�E����Fޝv�!G2��ځ$�]��KݎbŞ�W��G�Tyc�H<,���Z$�wI���H럿������1P+/@NOh��cL�b��)�O��A�^�}�~�3�Q,\�[�����9��"� S��P�nry�!-�u�N��XF>ڱ��7(Ť�%J���{˰(��m�AJ�A@��;���%FI�	�D�S:$�FZ��������~|�����^ǅÌ�ε�u�}�V�y�+��v�e�*Ơ�E�}���Ch�
��#��v×/=�PK�f��5��C�����[������_�������y��r��rrY��v�Jgh���)��(��ܛ��N����Y���x�|��s��/zeA���VL��6`�ڋ�^���S�t.����r��>v���]��K�'����d;LWTWe�A�#�u��ϙ�M��2��F�¾��z��7>����+�)ǒ����{��['�N0 �t,��� u'�A�)%�a�\��(7n�7�aƃ��¢ ~��ڦ�p���`!����|��  I�;.��"�|.5 �����'�����ɸ#YF�����]vE�	{�x�����]���R����{� շF1�k���YB\"�)�7hY�������1+g�iCF�ki��j��
{v|������"HxP�X9E���I֕��~x���P�{�(yP�����AF�~��4!���9at��)�ӯg"jf8IDܤՏ�s�\^]� VO���=��~a%��z��ݪ}G�&��,�	������
9�Ν��+-�r��t����{�8��d���屼��8��3�4"�G��j�K5���5��FHD}� �o}�+�$��9��8;��73;�k߀���a�)�#5�鉿���8"BII	3���5���T��O�źY>+�䮔">�C���A@�_Ι�|�A���K2��!��O.��P��+Z�O�4��D���8�ԣ$5������N��|9;7~��"���I�]���y�����Qizݖ����~6���*�yo^^l3�4�f�ٖ��4kV��ܜ�9@C/�_:�����s��lc��9�{���%�R��432�f�;v@v�+� �s�+���b$1�Hr�q��ڀ���v�O~J� ��c.�4�G#��u/����R'	��Z��Ԡ���S�6u��h���g��eВ�<��/h�R�_��������9ڻ����9��謄�y�a-��ௗ���o�+��
�hEت���-x tA<I%��`�������
�� %��}���N���yuN�Z[^�e�.c�G?���J%)m�R� ǿ,n�`l��X4ӟD�b�f\Q��G@;�F�W�4�S͓����](��dOJ��1��*a�%�"��V;��pgi����I����?bL��N`Y���fd�XA�D�Z��}�(w졜�#�	,;��dr^��F]�,�7 0rvG&	��p/���F��V\�YNsk2�� ��s�9"K��L�4Do��Wc��������r��p5��,�:~@s�㲑f9C��c���Q�j$�w��4��%bJ�О����W��>'?�1���p�N�q>ܕ��x��{Yn%�-#�}����Q�rni���j|Vdu=�XU�-�#�b�+`@�T 7��z�u�% ��~$}�܌��"�����&�C����*E�x~�uo�{�ξީ���6]e�W���Y���]A�8}Ӊq��6Ru�mp��[d���8� �pM!w���ru��"v��7��k��Vn"�}���]h�x��t�������^��B��p�{�c�
%�9���i�����qiI׏0!����Z�g��q��~Qm�a�6� �h�aq��0��%a�kv��4���4*��:/�[ovS\	̾�)߮a��0�Э�H:G��d0W�[��T��m���[G�kNNs�((`<���l�3b,�E^��3�*Q� JW�=�����U4c��.�!����CmI�r���{���d�P��O]V�[껾�3 kuM���ՕZ�`�=��'��'h�v����A~�@z�k@=�`������j�� ��<|����8����B�������b�`r�:9��,g���	#�z�J�ܥ�M�_U��+���&��8�U.-"	�E'&���L���� K.�?,?s5����^H�V@Q]�M0Q��#S�sR�Q�����plЉ����s�b-E�X~įn�НJ#������<]?��4�"�/���Ze��H��!4m���������L��0]����B]�ziw�gJ9����ej�S�pp	~@��j�X�sm�!n,����N૾��rX�A�n��F!�I���:�R�K��'�y՟����b�4|���os�q�o-���� �z4��۲8s���ܿ�� ����q�w����� ����A6����׹Xx-;���|��[��,܋��Y���G	�o��ݩ����qZϰO��{�Ø����|�ކ�J���ͫ��1 ػ�Y�w�j`$��1��[X��0&FXc���^�q�\?q�X
�����wB_TS���(��Dt|�V�'�|~�!�V� ʵIe�w��X��)�L=�͖W�����@̥�h���eN4<'� E� ���#�#Y�y��Qz>
sI�Al�����<�����y��+-�Vʯ�3(_��+~g.������.:�t��;��0�p��k���ay�"�,����
��|�G��.���˔ʖ�l���T���Rm����o(4g�jT譮��?����MzYUd0��>�|ou��vDY��D�2�*��TF-%9�)ӳ����O/�=?ߨ�	�ݛI��)�{�TE��"�wJh�+��@S_���e�;ӥă$��<�﹞U`|�J���k�P�QGo~�����U�S��&F�o;�aK�gFqZ�v�# O�	���O��8��RT�y��:PC<q�(�C��9Q��ݶ��`����?��9���f4"�/;�6J��|�.���i�e(�vG�.+���f��#��D�=H�?���������3AX	2�Kן?�G��bG%Hާ� UɁ�^�nr��H��r|7����N�<���i�6�ܒ���f ���t�Rz=�Ȟ��v5���.E����f<<�P[���2,��swH��*)iQ��{B?
��)���![�Y� SeT�Oݙ�l���r��+���Q������$J�q�ڣ<\:`��ls��"�,UXf�fURb��V����e1��P�,gP��L-��v�,2�G>Z�~T?���W� 
��s�>V���P�Z��c��lS?�4 &�\���n+���|O���d�����aY�� �Mq)��^/~�,	�h�v_��J�3�uA������7w"�:�J����@F�l�fh�xz_���P执�A�ֱ`Z��A�ꢠ�;|g�ǋ��t"3��ߛNh���L���cs����݀E�媶��� ��a���7/��=8��#J�o�������F�^�� � �۶e����� YYZ4ܼh���a�p��nv���a҃�p���Vq�P��%μ�	�/M,B/�-"�pJ�r�&1[���r-,�,�v�b�d]1�݊�b��Qj��T��B��q~	k��������C�۵�W�E�]c�]��<�]�Tr��Ę6�D�M�$*�J�ޜ�?��"I���}�u��@�y����O�
|��y�v����a)֥ff�S:�����i����:�u��:�-ZFQy�2(��ج�*a�`2�s\�8�-��-߬L����ba�����9I����P%i�:b�#��"��IL(�#�&]�{!㯶>��dt�\�㙵��
Sf��X��\]= �YB�k��U5���R��/r��[Xt��vy~	>!j���bG�K]��e�C5xy�n[�4�����w%/�v.pkZ���Z�g��Z@����Y����0��#�/�m�5�{�c���U����� �ہ���q�bŴ!�Cip�ZA����6+�6�.�1�n�=����o2����5�&$X��O)�r��[�Rx�2��|=��#�V�䘃�~Mn�?��f��F$ �B�c�
+*�Sd�U�1/�F^��A��U�Y��sob�k^%to����\�]O���6��^j���r�ݖ
�}-���O�Q:�u	�r?�
��M��iC9/�+�^��L�<Ġ��Q�(9���jO~�B%�k�4�5���SpFkT���[���bPp�ĈZK�����l�,ș!�+�B�� ��*;e&�S8����p��rY��;�	���P��hLtt�����Yה������b��Ww�9I�5A�>!�Js���)'/&zZ�%���kg �sz�]�fjZV�\�'������އzl%ᢙ&.��[\t�o9���e�t�a$���P�(:��WQ�\s)0��άc��0N���1��ೞ�S���;B�շ�9d6}���U��������x��<�X��r����c�s�iGۉ�'�����л�YM��1����Y�D&��B'�C �o�5`ɻ6!���ǁD&��{2���
�\��e.Ҥ�D�^h�����v�f�T��w9QN��1i�}����;ӏ����&�"֙�+OU�x����&7 �����.��X�ו��:���N�������&:�m�=6�������b�"Ù�>1(UCG���n�q��f��mg���z��`��!��&���^^_�$7'<WLv]�n����� ��6@�Rk����-��3�/_��"q+ -N��!S:@˿���	��=VVI�p\
;4�|���y����6�ѿa�� ����R��^�HG���X��C����x�%)/L�"w�OiH��<Y���Ԯ�	Nk>��xx�p�~і����^.k>�O�um��w�ڜQL�yRt��2��}G����.Q�Ϯ�~���g�umN���+�r���8b�+3��w��(�Z�����eb멅��85yd���]p@��M�dtf�c��.�p���/�m܄,�<��>H �W�RD�,��]��6��d!���Ò���ΙJ�S�O���_�o�!6�y�[�5��/i��e�m}t�YH��#F�8��Qa��Z��SN<�0u�r�r�Q�AF�K��i3�3�N:s�.-�b`��-��Wl�bw�헞�Vί��b�X(A����ǳ�n��N�.� �@,�vG}N ����=w��t(�r�� ��n0S��T)���J���d>I��1<A�X���8F�Q�����D�\{,0���L>�c��^Y���3���yUĴرb��Y׈��	��X�U1��[�8�ق(��
������1/�ۉ�%!֥k!3��Dn�+�����D΀m#H ������*&Q�RŐs�F�껓Ʋ����F����Kˮ�I�����uͤ�_> =5Ӯq�|2P���@���ak9��כ��]�;X֗�1��
m�����	�TP��)"h5�?���EJo*Hb���n�|�*[$仨;��
��?���Qad(��(A��0��0���e��]��)믗Iӎ�t�����Ut�����z$4��)�ʛX�:qp����ӌ�s��Gl��ʰ���#�85��h�e'B������*50�4k���o#�+��H�
��Q#!�����_(C�a��L )�M�����!~%N�XꌿO�*Ղ��ܗr<�����{����I���?��[�qr
��4T���G'�q"�:I�x�!ͪMI'�:�#��2B]���4��g�V��U�*����P�(p5�I�Of�Z\���r��`���a�]Q�y�w�1��Jd��wx����{~�1@���TY�Z^I�#G'J�~Jb���������m�1�I��$hjH''��S��N��Sɸ����R9_�7���c��=Њ�Q�<��.���Ć���D��NX���������q�bx���n�Sz�;�ZfջS�D��}��BP�2�ķ�%�&�t(\/�괮[�t��P3djeC���ҩ�y��gg!x[�y9���9WRf_��4t�^c"u?2:���#{�׾�q�q�4������ɺ��s��o�A���1�j1f�e����d	g1��9�z��!edyJ�X.t��4w;�)�p>jX���Q�������إ���w��s(73*�bU~�CϤ]D����#)uI9G��#�(�Սb&�C��C�߸�ê�؀�v�sI��MD�\9� ɬ�"��?���}��qص����eOE�&X�#�?���˞}��ZU��As~!Γ��;]���Խfk��)�=$_���I~F��C%��~(�/>���17��YV�Z��id��$�q�^�Z���}�#R��z�g!�QͰ�<��iC��[(x�s��㘭�B��;�<�z���2B���L�$m)���j)�Jf�Վ��ǀh�p��[a410:;~��#0��'(c���RJ��������w��<�U(+�˧s����!��HnZ�VD���Ed~q.W;K�M�T}Q,���������v��;����bU�X��l�b�	��Cο�X_��%�L��;>r�Y^\<�$��op���?��eR�H��v�X�?�`Pph%@7��s��E}3a�iH ��|��(�1}nҍiv�!���d����;�\�~Oi�J�na��I�h��7��i �!vy���^���ލ�r5�T����\q@0��] @�^M�W�J�U^�H��쥺Eb��:��Ȅ�~��O�ƃ���^��5��L��S$I��у�>�*��kT-�~��-"\\���D����ːbGs}���ǉ'ňyD���	 ��b���X�2Cb��9�"��_K%�{�<���C_ �T��!U��I���ǆ#��?�2J�)����k�J���	����"��)V=���mj�~(6�Eu���� DH�L�x �����w3��o�p�<*/i����T��\%�Fڅ��5��U\*eٯIX�~�yIݏ���s������������{5`�l*9��
�,o ��v���od�������r(�����?�A1zk�7>gDHOh�wQ����p{� �r�SfgGeDx��*P��Up;�^��^�V�]3�و�rv�?�f�L��9nK96t�Z�,0��oMr��Ƿ��Qd	���H'��%43V�DE���ys��0����$&��E���E����~�q�1�W���L�|���E%!�%��J��ְ�S���5�C�=��aM�4(~#��-��'��[���+�[�����6m� �����D,���ﱸG�0.�+�-q7��q�olb��rtݡ\+y���7��y�#�����q��'�����Ȁc܏�B}7~u�8n�\4qbA����-+�x���N��i�Mv!���La����ªS4�iYq=���J�4���I �FdKd�}!��c3����������Y�A�����Rb6�T�\i�b������ `�R�ַ��[E���)w&[;�� ���Q?�p�9�����Գ����_�=�������ZFS>F=�G0�8��\/Sӄjq;-����3�r"����gǳc���Q_)wv��Y�jm���p�����(��z
"�l9�!Q/�~n�c���.&�:�`�d��y����x��4�fWRN�}6Gַor<~��6�*��x�j0p]/?ev����C�<�'�8�V�A'�:������j�����;�!�����_������!�Xҕ�g�]t!��4Ag�mO�����Cli��8Խ¢�llV�G����$�����P���yt�d�yZ�HM���k�s�ojٞ�j7�z�8��_�uޓJ��&��[�ˬq" ��G����.�'%� B�ZQ���с-�Ah�\�$,I$j��5P�:y�8�pȥ2�,��r�^�f	 �W������4�^���o�ƒa�&����5[l�HߤV]�S2z��;�?�E��72��YP��n'NR�	�|���Y &1�g�`�����|̏��K�ș�H��| �Z�jv���b�g�q<�J�	1�����8ET̿�#)o��b,Zwu��',����d���mo&��R ����̧5L�5,�����?㞗���_V抠#i��"�ϑWbe[��$�s�?Ǯp��R�7!��LH�-K9D�Xd�m>=+���ƿ��\@�>�ڦK�'=@h�V��M6A�p �"���H��4�x�D�y�=
���D�'��u��*����(�R���p.�Q}x���>@�Д��Al�l=\�3����`)����G+~�j���ɿ�J��t�R)_v�,�4�n�Z�~ERg�to<7��a3���B+��6%�{��$�*W��K��Uz�#�^\���3���ґ]�"�E*	͘;����t�>�^��Jy�P&�]��������]�����<��9�� ��� �Z4��\�0u�|���)�P����Mѧ1��=죗���_;�݆7�^�Q�E�jP:�<��a]v:p�r_T� 5X������R�=[��uUÖ��6\r�K+�;T��
��/�ؐK�pj���q
�/�2{��D���$P�����L��LN#���b9@©gW�譹c�y��8�ɲ5�jb���<�Q�撸�%��p�� $�>3�@��]h���yi
��B
DA7,S_�,e�ȀVZ��gh���rF�̡�uщ��%����ݣ#��ZJ3"*����66V�1CdZ���Յ�U'��odte/U�E5'��S�9� �ac��gimE��f�zn���N�q�]XH�"+�*�D;�R��*Pmq���1�����+_ͭf�r����9��Y)�R�wÔ�ؖt�� ������`���j܄ޖ؈; B��`��:�i^�q�O��OT��5%���s�W��G駲� �O��v�Nai�0-U���7P`]�AS�A�S�O,Eu�e���-�	�2�iK�Z�IGiő�3<�1���v�x&`�,ќ:�3���c9�_��)�����S2��  |N	߇�� Jڨ���D���Wvn����H�$���>Ǩ��Ƭ�ٖx��論;��ܦF��g*w�z�#Y�L�5|��������e4�et�U��U�����!�'�R޻��u��.z�,%<s�]ˉ%���舁�J�<�8��,�������cAY(��,�~(�1�E�P������56�"��ϥ��������CR�]��x��-�Q�$�Pҗ�����7��S��|��\��O.?Ha�������ko���Ɍ*�ɬ�M�;�:��|��s�c����l�B`����Y�T f���{��T�����*�'3�*A�71�?ZHh�����a�3:�b��J�OU
�G��#���w#����ەS��:�_�#��/f0B���=�B�A�����h ��D;ƌ�NN,2�]�y�������N��$�z�2����U�!��F����b�dL��K��Jф�MϮ,z9�s?���
���dY:&à��P!������ڈh���)m�uh�I;80�Z��`� Al4���]�C��a$Q(H�(���g�j��3��o�2Kش����o�T1(	)�ۊ�(CY!�v4N�����s�Z�a���9�ẁ#y6��3s�.�z���*�3��20����D-XyB�����G�76�qE)@iy��8��8C�P�sE	��!��A�8XdA�Mj���:���aЖI�F,�PM�ޔ�9���ҵ�Kz�����/���d
�N�?������珗!��
���#J��_������q��o��~de
��>t5kGs$��Vjo�k ��Jd���ƣ�,뛁��~�M%(��rJ8�X1�.v��c�����c����sCr�ML�RY�N���׼��B�����Kѽ�����,}�� Z�S;����pQ�J�6F>)�p��?v@�wW'�	,����C_�zzz1�Ro������q�%�e����0Ҙl���c��X��F]ʰ���|V��xi*aC�Lq��{|����xjآ�i���(+P�{sл "A�gMFx^�xMF�x����x���Hf��$�JY�(����%v	��a'��AI*�U�<cy���VL	���gfe�51Ɂ1�muÏ�«�����`N��K�^���UF���d����k ���D��Ś��H��A���|���.Bp2AS ��Vnt��p�a���_��ŕ���*Mn�)��U�Pr�h��۷�C^�-���Na��Ӄj1kx�bkm}�ǮYD�H�z�al�&���Ԫr9�*���}^qw7V}�*�
�ʦ�J���b�&�Y��KGL�`,T7���Q��
؅X�*ϣ٧�"і�@+��ߙ�9�1 �B1+ˊ'kͫu��O^�H�ǓGn'uzg��P\���(܆U�|k�!��ɢW���}�i/���\�*�+��tD���W��k�V\\O�l��pN�6����M���3
n�#��S�O4��U�
GF2?UH�bA����_1���g[b�i�e�B���r��ȫ�{di!��k�vժ��!jp.bMD�&�z���B#niXDH_��9R�'�[3k�H�{,�y,Թ벟�	�4;�#�1E\�UNçJBwk&_^^�kⰲ��M��~��a�O��,��������7/�}o&`�.�P�P�����0��Ĝu�]?p�M�D|j{ij���0Z� p(4���̌�R��O4��C�>|ȻJ������2yb�2���ڝ7r�9<�>oks��4��̏/�46��y�A�����'}P� ��3��w�[����d����9X4�������G�p�>;"��c�t�.����'7�������'��9RP։���=?,���^�4ާԉk�2���+K��З���,�����2���g �D	S�������$�<J�XXY������_�Y� ٰMG}xpՐ�(�p���{�sz2��L�o	w�טy�B��}�ׄ���˷��k�y���zN�%<������n&ț/zps5�� z ��T�۞�����t�'\Zqx�/�da�.j�>̋���j����!~�����"!))���#Dct�������0�����''�oֽ����B��6OD\�n��r|!�!�f��<��8��'���De��+b�|w��jP�݀�[|!�����9շg��o/@�zi����"�C�֮g5�W� �������t�5$�mO%�7��ٟ�u?�T3���j���x���䓆�;��Kl]�+G^̰�(I�/k<4�$��kj��7o2�N"xFܚ�Wx�,���Y�x渷�!���k��@�,�X���w��	�]�/��xC� c�� �rs ��-��]�V$tp�2ċ���2v�3ο[��1$�hD��x,�.�����{���sj�h���~nڭ��4"�;��M�.jh3��A~�8V�:"��0��'��ڨ7,��=�e���ķ����p��t]�oN�%1I�(�?<�Wc0O�+�(~f)V]�>k�n}��mq�# ���̈��*P�h�0 n�l�	�ytU��Z�;�r����f���b����U�Y��]��̷R��e��:T��|�p0��S!�f�n�Y��1J�n��;�|24�y�6�U��c�y�5P�|+s��d.�;�auV����o�3&4���Û��+�:�	y��Ps��К��2չ�]��DYlZ��c�8��p��$���	�<�'�����m��,q��7Q	\�Y����nܥ����B�bM��[I�E0��А�5��f��T��1�ܶ'�25�7{w�!I\%+L'B�uQ!��g=15a�Z@��մ-
�@�R�,�o����ON���W#,˘��r�4Ù����jas}5��_h���Ŕث�:������o��q��WR�zn��~�jSYO~�v�$O�	0 ��?�������wB����t�͖3��@�hG߿;HU���Z"� �}����j7�gO��)m� <`.^p��
��0K2�zr����z�.O" �X�a�$t}>J<��Rg( �ц?2�8n�{����k �z	��&�Tp�-z��4�ɺ.`2ſNZ���Q���5���	�3:4�ε4e{U�Z���]��?��U{�����ƨ����r��8���F'ʦ���?&��U�%�^�)�l�(M֏�l�RzE
�Rt!��i�4��F��}�:���g�����3�[���*?8D&U��
��	���P����{^pieI�,_���bG%����������*W5򤴇��%e`�����bk�
x��]���ԕ�}Ο�,�C��g��h�Y�9<�ì��E�y�u�%���_ɹԙ�T)z��~`4l��5;��Mk�����KBL�$
�F�:�tٓ� �����Q� ��ҏ�`�=�rM��O~GvL�0�h����"�,Iv�U��Rn%H�4}X@���}_7��׶O؈��NQ3z��^re��FUד�;g���.a�dI��U�-��$3��$��#Ԕ>s1jr`�("س�f��ӭ���^��Z�ԩ�klǕ�{,�"�K-�E]%��Ts��w>c�GK�/�o�hP�X?I���$�g[Q@���n��r�X:��t�*�89�P��F
�C���ۇ#��x�hW^����Κ�u���S��Ks׹�����v�pٱH�Kӕ�F/yS�n��2�a�ۆZ�F��Em�b%����I\(���)p�}~���f�êo�ݾܦY �>�x�u��G���:ꑯ���P����sJY/~:�PUlT�e�rhL��x�[��q�|�z_g�_�.�?.����
D�6[�]�'�d"4,�Cc�+Y"e�#\?~�)����3�r������n��>�լԇz2+d_�3W͞�(��rD��c���"aw+�ی>���+�-�(ݲ���}��3ϟ'�:xۗ�"���Յd@�;v�L[f�����&�������H����i�;8 ��'4hI�p���|�#Tc�������b����Zlؒ��bU~��L���esa�-~RGO�~T��[�=�[;�4n��P�T.��-�ծ�Ӟ-e����D�,z=���HI0�a�1�u6Kp�p2�uI�3w]��[�IL�5�#��<�ҥ��+6lQ����y/x��o�<&�,:]k��qu�f1\ڥ���Q�ӯs)�����3�o"�K��F�j�U��b"�X�4��~�r��щ�iK|�z{����?��̚�Jl����}�U������@��z�rH(:�׷+�r�����X��kS��א„�T��
�j�4��W���-.��1/�>0~&�}�HE�x�,�a��Y���ON���(Fx����gse*3L�0���N��Ջ���DM�[���`����ẖ�W��\Oŋ�$��?�oy�{Di#�I�X��RBć痾[d{M��7�!��Ԥ�O��t�@���ח�����M R{��x�N?Q�M�:��Er[��0$��|�!	�X�
�,�6K11��PÂo(�)u~{3�PwO=�A$���`y)!�����E��y�)1e��ԯ!���n-��~��2�R<�$�%w�r���Z<xNr��؄�_}<�ZKM����Nyh���s�'éA�Q���$���x�%Aj�t�N�i��;���m�\J��9y�8�UX�t|�'���4��I���x��}�ç����q�'y�]Tj����j��.<�^,��	�ړm���?�l��2YCG� �3���x��7l�Mʷ�Q�&N�!�n�΁{y��+�<�X����}�x�I�ė��p�<M�?��2���H,�G�%�D��[5�96}���l�iv������M�~3�x8]4�1m�Pnf�,56B%j�R
�%�vb�e����COOK�O�'3:���2�b���?��������a>1�E�&B�^h~��EJy�d���u9j!ot<U��rJd||*�숤-ƴ�+�.�~�9����Sw�k�y��y�K����G�%��Q�� B��:&x� �b����\����W<J�cj�e$�2�DD�S�aiN.R����_%c�I�)f���36E�wV]�'D}k�M�J���6[�@�9|8W͎�J�GݟK�=fP��W̗-]�b�LG?�!���\���l�}g1k9�����x�3 �I�l�����?��y��f���$�U�o�;!���ש�����3��0�+�SY���.ޞ�hpX|F��K�l�����F�AXA=��||�cV�Z�" uM�yR�55���N�&r��CQ7���s�
0L�mI屳���$Xz����aG�F�7�[��_�qUG=�^���)z@�UzBt�i(,[Oi�M�����{EW���g-�?�~�hx���w�վ���� �mk�urL�S����~��.-n�!0͚#���:B�"��9�A���VE�g��k-O�!�2��q�ڹ�A��y��{ħ�S�h���y?��(���R�;1	�t���"s���54ZU�,ltFD�.�k�y�;�bO.�LI�@�#"*XP�L=����g�ps��F����:�:g������OjF�Fr_�ޖ�/'������C����uޢ~��XP���N��*A
���Nl��+���������?k(�����n��(�[Ԅ����j:�gN�:�M4���~޶����Kܢ�p��L�<fu��Sٰ��՘A\�֑q��H�&�ȇ[��zʍ��,�I���u�3�:�����qQ��~��+*B��υ��mЊ����Q�k1_��]��~yEZ6
Y�_��T�@U�||zE�$2U���(�۶��u�a�i}-�Yg_{�p�64v/��������y�2i�?��]���X��e<^�;��������ߨUZ��TlX�U�R!�����v7�ݥ�d��%��wv�y�f�Z����jGG���	U�߼�=�A���
�ur�$�\��_��/?�ou������d�k ��3��0��_<؍����,�z ���yЙ��i�: }��<#���RRh?�?��w/>��Z˼�CO�#(:���}pu������6�����ĜJ���Wra/.܃�7i�{�
�y�%`w�W���Ґ7�+�A��}�Ń%�#���
Pe,���z.�ܙ���f�{��	Nb��j�Z������Zd3�4��]%���:�I��G�/0f�K��D�gC#?�0;�DԷ�7�Y�n��8^7E�}Ȑ�C�7����+:�5{����������ga�C�$ ��NّJ��_�H��`�g��&�>G��@׽,��]�ԩ'��N�:콳��"�^?m�
>�o��\�GF��q�u��*�#gp���JQ�Ó툌^����T��b��ABt8�n�s�,YrFf#*��M���з>?7T���W�ު{�,�w@�n�}���oA�=K��j�� 3�����8X6��z��� �5'� �Fz�сX��,Ѳ?[;�1�����Z1�7����2��_+���v��S��F�����NJ���y�T(�V� S��.e�?doVT#N��~��%�d����_�B8�tƱ��=:����x܉��l��}۬^�����L��,��7��EiA��]��kB���@���l���t�6�o"U�'xpZ)�� �񼽀�{x}������(:1�;q^I���<-3�ۆgx_+�)#��/�� #-��ދ�_?�vn�ͷ%��N塗�;s���e��Q�&r�>k���Gޒ3%��ۦ���	Uc^����Y�xc�1ѻ�$5�)����0�#v-P�i)�E]�tWOg���JĲ�<�;���P�]��Pr۪.;���2�ik�Z����M�g)E�����r>��@#�d邡���iU�}5�{��'����ib��՜���R\"WS?��ů��@��ή�Ȼ���e#]���Ӕb��S^8��L>�G���%�}�8�4��{1	�K�i�
�Φ%w�����J�[��F���%�����_�CGAB��t�;P������t�a��V9)���K�F�/��� "�i�7+�`2� ֵ)	i��w�P��h)ds8q@�K���v�&<̆��R�r����<=O�>���t���*�����;���8�^1��888�5��Z�?�`��,���#��޳��6�鐼��g�83�Ы��:����=�Q2�J�B��c�L�T��F&���.�����d���TD��7�?���LSO�qxi��%������B6��h������hx�M��o�C�燶(���P"��}��W�T����+��C�OAAe��s��<�)$0h3x_oO�A�H��z_�Ұ���O�!>���
~"w���E��?�������~�0��O�aλb���D���[�K�,"|�~�u��K�
�� ���8z��������Ub��;��L�%G6����\�!��I5��7���;GM3���]R ��ѻS�W�}f�5q�l�T��"�V�ćVȔ%�
�߉�����JX嶹�϶�|�A񗠛�G�U�
��&���cѥW,���AP<���$>dbM�U��Koa/��}�����X�v�
�{m���W%lt���
Ɠ0���[pއ~~����g2;z��=fո��y���;L��k����M�,'!J��	�_��� ?{y��UxۜIX����w:�*��jv��9]]EfI1Tď*�?>�m�����~���|��	IO�l�&N|�'��Cm�m������,��>p���B1-GD��+LL�5l�u�����{�UU��Z9u684�'�N)��䶟�،4��vɶ����3��Tfj�8z9��gWOO�H|#��c��6�܎��Nk��#aH�J_�˝�Fm�'hal2C��&��ق�ſ46F�#0M����O�U�e�WWG�x�,��?<}e@T]�6J)R��"�H���H�4���Hא��1�HJJ����w��y��af�Y{���]���ߪl����l�;�t�Gś&������-�c�N���x]����q��Cӽx���mDBmi��wP'�3��~#���6�y��[[B�o7
j�K)l�
�p$+j9Ҵ��	l2�E�+#ӥ,�;�p�|�Y����Osk���{*�knj������uV��X%���EPF?dï���a�nڷ�4���*��lB�p�(��]Ycss�BO7�>s����AF1�Y5�������9HJ��ճj''�`S�5w�y���ŋ���T�����������i���S)�ٜ���vG����_Ϝʴ�m�,R>�~3���I��G�wW(&'e���a��4L7�"��{D�#*;�
P��=kN<���1�gM'��J��Qĵ�la�: ��!�*z��P���~A�bs��g�/>6���l��`�(��������
_MQ �#�2���?ufo/FlD��jDq̟�K�q};���gR96e	�&����c�f<>����9���j1�bdAhqtUW��xW[���y�,��P萷ȏ���Vꠘ�m&�oϐ,��:s����k�����k :����O���Ḱ�%i��Ҽ9ӥ�&��!����u�#n�Y��&W)��0�8��Al*�;9&xQ�֪B�E2X��g�Uq���9����@��� �=��B���jz���7��O��`�= ;1W��H��#_sX���"V%�aNfL�[\^�����I �2�K�����o�~AK�W���UY#�	�岥�o#� �G�kVR_����(�6�o.++��'��hOB�l k���V���E�Y/�Ë,�:&mк�|�hA[����z�^���ۘZ"N�.r���b�<�`i�3�F��\�=8�q�vbL�H���/�yMm��Cosa�֓���G�)ҽr-��BV����=�p�	�d�	�)k�����38����).���Q[�ÿp��M�1z�$��b\�<����8ۄ��BnH�n�1ϧ��0 (Z��o�x	�5�G��^ONOK0����MM�����LWQ~��WXOO���H����'��}�Կ�Y+��a+ӱ�wS��s��(�]�aN�jg�p^e̸ ��<<a�<f�:>�=���E�>h���$ri?����/H�XtΐM��]������=�M�X���+B����B�06P.Ç�*�%*����������Z���2��5{�[AC�?�!�5{�m=�*J�[*��r`-}����sBw)����1�v�����d�����闱���w~���Xt�	>F�H���C��#�������"��f�ySnz=׼D�E���Y��!�P��kb��ȝᣮ6~�'n��gR�t�B-��"��C�T�|YU0% �<�������'�����Bf��O��)#��������^�ә{;�~�|�j;��,�W�|L)��J�vA�$r��3�$d�Zu�{�w��F��_���`{{���Κ�k>� �/����C	l
��(4�X
��ۋ%m��$�o�-1	I����|I��נW�v@�@�ŗ5_y.>�9�����2@5�c���J��Q�.�*�t;0Ss�<�1۶�h9o]�R��*NA].��-���VP�K��7β*����e5�b[�(��^�S�JxK��
�?��Dz���@z�@3����]&C�mt����� �+�/���팀�X�J�1���z�y��r�P >@S�7	�}=�6P@k�R�E�����M��{��G\'� f1��ص�T�Q6�*��_	i�����,�U���}��u��|��{;+N�Emx̱`�'m|�
�� ��?�.���0&/[�D,�<6:꟞NE�%J��m\�� � ��PE;�0Sl
��+��':#�`S3d�WgFI����P�T8R7:f��������V|���]�a��l���/*�O(�#5"@܍�K�0a��F��[�*Ro����%u6�5��a3r���Sw�l_��<=�ˉ	���
J�����j���~�.B�5�p��g!>pʠ�m:\�
���X�i�*;�ؗ���Č���э@/������2l��I�d�d�W0�i��KG����c+��}d��φ���FK��,]�:��Wlgw�pP�I<�?���'n����)���6!�zG4�A�����m�cJ탄��3E|�z�����BU�c�l�Y������Px����_m���zlp�w<��S�T%f�Df�?)�Z�5�o>����vx����Lݜ�٘l~n�{P�����P*�T5Fh5���S,*�_��$P��>�k�n�!M ���o(�Q��)�$�
��ΐ\�fI���|í�jS
�b��4W�g%`Q�����fUE�Kdr�[��*ΫL�=)�?�o�����x�"
9L���PkN׾Ԩ�Xk|�ʠω��Ə?��M$���]��$5��M�6A����Z�Pq|ͣ�-{r(+C�F\�Sk`�ǲ�X&s���2G~���l�"�w�ާw~oq��8��#&��f�;��f�W�s#r̼����t�|�H�j����_�h�R�W���"��!�.�E-�e��*�B���@���ou��o��[��ei�g	�@R��F��3�($��ջ���)M}óm��w��P䞌�`�Ȟ��������Y��-�2��EO�\��`�A�����B}�II~��80B7�T��h�T��R�i�Gt$��W�"Ǵ�Ϟݴͫ�D�-I��<J�v�W�:�a�`e3�N	���Ģ~�FKc��C�za��m�,�2�tM䔄��%,c�n�s�>ȡZ	U�q�V����|��_�R�4n3����}�7${CV�s�ӈ�d�߇�*?�_e���RӶe*v>���7V�㥍��pp�Q�i�̗���if>

Z�;ܙE�7����
�[��E�.���Q 
a������Xxsc,�a��A��b�?¯��{��z�bL���~���x��8�W��޶�R��n-wV�n��^ً�W�����ѽ
�[�2��^����yI{���)M�����o��O7����WY�-���e�p\^���[���x�L�a�..�57I�p�2���l������N����m����**�;��QL�����qQ�+M��T�<�h�$��!=�vO�un��Պ�B�9zjU� ���jt�TLgX�;���6����R��3���6��)_�$�_�����ωq��A����r$�Կ��'��Na�ެ�8A�AoO�C�x�B���Z4Y�ѧ���[Շ쀃y����kU8�QiHP܎w���'��i�-7��~Z�b��,���:ڡ[h[`�ڌ�������0�4y/�V�\�Z����by��ԟ���$Ȣ�/o�DD���(QD�~-���n���6�.�
qh��P����M6���	��[�to����p�o�X�����c��.�M=��%�A"�Y��$��;OR{��#�<'C"������^���Ŵ�̆�=A�}�dx��z��Jj͟QHړ!�,W��Z8GO5, =;hw�i�l��H3 ��d�9i��'9�������䃞H��i@��ݞ��k����t6+ȝ7
U��{sa$z���^�0�Y0�K`��=EIL7/&sc� C���a&�,:r���Di˙�$�5��ɜ��A���Py��ЇuA�(�Vڈl_gF�B 8�p=^�<�����ٚj��/	A?��0Np�n��q��2&��?����ي�n�Jا�\c_Km������ov�=�gǕ�bݎ�!=�b��ʻP��������$�sv����&L��V����'�<���0�/;�bFNxb#�|ߺlGę1�>�^���
�.K/LUF��Y��ʿ@3�����5��i�Y�J�����Kޭ��0�Ef|�|5Q��[�q؞m�y������1Q��'�o�3�ߙ=���Qcr��Hq	=���q�G�ҵ�����xV%"-&��?�_*?e\L识/�{2�͏�Ȣ��>ͽp_T���ff�b+�����W7վ����@6l8n�����Kᓽ�wF�ø}��H\�l�������1'9Lԕ��Y� '�y���W?R}nG��6;y��-'�R����'�}�Z8�q�W�=���3]p�pܹފ̠2�7�V7�Oj���5��35B���w�p�0e�v�ԥ�]�v)�M���D�i�|S���Y���M���:�A�w�F�1��Ԡ��u�`k��s��c�]H�Ha]B'��n �4���m�����l�E���y�{w����r�9�氟c�4��R��3�v �G��ոt�q����+-�/��K#S�KUU��a{fO�0�$�.�]���5z�h4�{S���L��Nɐ����oٟup�`���~�+^i��V̎Bp�Y����z֭���p�<�Ld�>$�UQ4dP�ϩ�����ba>�4������H$h<�������%���8�;�� ����~�(�������J�T��alK-:�G�si��Mk�'W0�4���7�^��O��>{g("ctxnM��-����+�aSA��º�2�B�}����y_���G��f�@�]�-]�|���Jܱ�,hm�~� ��RÃ��S���c�@w?%��j��9	��U���l��:�ʙ0��^޳�=�/KG]��o�V�4�O[}&�& A�O��J�!��	��w�"п�!;&�d v�c9�{<�p��wn�级CH��Q�Z��_�9��t�?��& ?��Cb���K�Z�� ����;7�� �c-�qA_/=\>^���"q8m�l����e�Ƭ!�$��>�W7'��a��i�P���`�+(Twlq
d�+���žc�9�U�/e� �M�$�8������L�/w�LfK�z ����0�;ߛ�ԽNN�6c�i(��ڨV�[@W����v�C:��v`��o�W0%-����F��R�M�� �<��v)�e�p�1��e�8�%��bl8dJ}R*R"�젩�}=͟^�g���#k2.�����t;����*��U��lg�cl�RĂ��\I�~��1�oW��,��
�M�����D|�&�qI�����ǲ�oQn�.�T(*�A��Bx��#�M	��l���.�)7�&��1ql��pO-w"F#Z	���=?�{�v[��-��w�������o��gQ�}	���CU8��0�ԨH�i�����*؋<7��N�p�h�GW����"K�ھ�H����\��{8�~7��P1�/�|3�C�d��Vvr�0-V��	|�Z?�\)\����4c9$~|�h,f¾�b�u��������O������Q�j<_�
��b��!�I�J��F�\ӹ��p��Xĸ8\,�gx��|�&��E������(��#�h[�ЧX3�S��I#�7�)F�%�fI��2����J�p�^�~Yjy�+�v���kK�R�	�&6B�l��'R�]w0�}�k님�.���j�������P��������%{���o����)��u��(�A����|x�J�\f��^F���d�u|X��S���@�O;;�e�����9�������ƆD�c0Q{�b�U$��x��� �EU����b�</ҫ���$�㋵�讂)�̊J]����C�yu�0mY��mfT���ܒ�����*�N��܂٠�;�'��ô���i��������
��7�ym�QF�(ڞ�@5կ�YE�G�m��0���:Z��&K�ӕ��I�_o]�ʹ��mO�g�m��Js*�MqIȇr�}��/��\�/�	,"	ʙ�H����}V�.���Ԛ� �����l�E���R2�Ǹ�99����tu�5�"KR���4�S�� ý�4^��M$��C鑀{��1�����hz���O��į,��4����1���w[�q/�Ո$�5�۴��[��Og���(�OnO�"���/��[r����j�2=)Cx\:��B��@-"�	q;șc�@L��(H�#UpjZi��=Z<E�l�er�
@\_F�>=�O�Yv=���,%X��m��h�ĂE�fNR?�MlJ��)���П'�8ew��{�����Zx �0kAMK�C(� �O4�ۊ�v�{6u���#q�����v��$ט������[�Pmo#Pr�o&끬���t12p�3�I�15��w&< }QK���K�TO��X�y2��w��N��kә#d�U]�Y���(�����$i�kB�5�_al��ܦ�L�����V�V�vx���F6JK�ϭ(Y�,#v%&�Y�͟uOy�G��]���d��"��b0��$���'�gU�i���]Ȭ!�|r*��DTDOl(X���x=��63�)��^m_�ڜ������I$��/Yl�6���0�BǮ�_3D�|،��"�W�pb�˷!���[���[:���A�7�4B�?�챳~� a9I��ED|���>��mF�T��$���<�Dq5�|�57���Ҩ5��K1���ͽQB��Oc�M���T����H��X��H�LUؾ��}���jR�X��C�X�w2��Vs$��"!���݊?^���p'�q�=�R5�7�\-$>�;��#��O�Nz���X�b-���`��J<C��7;e`SUb&��@X�D���y�j3�jEg�ߪY[N��
rI?!�MF�d�_�K+*=Q������rt�&51~�r�}�H�\K1�KA���·ů��yH��h�M�7��gs��5R����� ���d�J�T8N��]���g
z3��E	�_�����>l>l���80�����<]��k\�u~���^�y�&��O��
%���ǉ��� �*�A��#���߹�������}��l�SȾ `��>q~�f��{�F-� *: ��_��Jʚ�7�X��p:&�I(��0�d���x��!�A�E
����X[�����e�<˄8O�%pܪ0y���6GfL�l��9_�!����a�aw^�A���-%�W�`����3��Ow;�RWUEj��~����D�>I�G����S%	U,:"k��1�V�C��S�>��}þ�m��5�-��>q���b�밻��[�)��d�6Ԏ�@H#��W�RUɿ����B�������v����؆v����:���B�y%z��KU��0�����;x!��-<�{��9YY�	��v�-��̘�j�����*+�Z#�Md���|��u���@�O���F��X 	k���9�f���◁����������<_�GqF�Nx ٰ���`��S�G*���3����z����Q����LΦ\)�YB�u�EE@k��S�ď��DZ	D��Pu��tR��K�����h��hI��`c����s���+D��Mߦ^�����:&�?X~�c�[K��"?}7�M�/<��^j�[�Oi:ڌ$���
�� ӟ0�PD)��Q4����Wpm�|��ȏR�R_��;S3�ůT�PZ!��Q�����i��)Qj*�j�}���v���c�O��=Q���B����=MQoM����"k5J��p&���,�������6���Z�Ue`z�,�����%Isn���y̯�4B��Q������C�+��5S�^�g�'�s�N�6��8���rr����2zݦ8��ay��gv<(���h0,�@S=�ˁ��#��ӀB���N����>g��|���Yl�Td�'�ڳҷ5��7�6��e�R�S�wc�8��vt��ra�!��;T�u�$�����Χ������v�ֲ4�3�wE�_y}�������)�D�@�AAQx���[�4�,=?�.��0^�|����7tM�A�F'�h�� $!���*P3����h���O�/�kh��OM��sa���wOx~�K!��m�pQ�L�菺V���U!�;�kAǹ�ߐb���g�#aUVt�8u���8���: ۛն���={ԣ��(�裆_$� �c1W�Q�jr����wǁc��g~�㖦��Q����ۍ��Y�Rl�Z�`ZD�i��?�M���16�Aܵ'�G�Et`�#f:�-�s����~ME�l2cTB�D���;�sk�2�����巨���,�Z��U���Z�֓kmg�E�O���,�E�z����.�$"�F06���ʁ��|�nGu��z9���)��cp���@��j�?F����r��r*�(��D'k��G�5�j_��ig=Nt_m/4�z���_ډI��FWL��ׁ��"W��+�;�����f��I/v��eNղ��������b��!DM+�e�mr?� ̩J9m�x⳰+�g��ݢ2<�k4ֵ�� ��?�Qu�ź3�ƕV�҈m��j�*PbN�TrC9uck=<H�msm�)��C���������l�o~�|���ȸ����QᜇY��
�]�1���K�O+����\%u�V��u���!,�T����� ���)9�^�p�#���%��`���׿�]Z}��(h"l2RR�,1H�tDDD��Ԝx���ga8�:�����rɱ�ʮ�@}�nl��O�/�FekTVߟ'.���-��ʟr��&��yo���k�ˋS��F�YK#����P�t��a�
���i��ɺ��l.\��d���*J��=1������/��aM���ks�DY[���Vx~�]�}_�p~ ;��l�gM�?3�5(��PHRB�ި�=ó�m퐥�%��N/��M[)���U�۴Ƕ�<��dYq�?"m*/��`	�E��ۨZ��;u�wwn3#��#�:@ ����$i7A�{o7I�� ~�^����"�?8~{M�ɦ�A��a��Q0�����}��)��=?/�ή.+Q
�g�sk��v�����"F� ���J'A:vOI��ꖳ�.\A>q[���Ȝ�7��,b���(O<�!��>�.�~�j�X����R��^9J}gz i���ɒ����� ��yd6�Җ�1|Vm�~mɹ����K�����3�u�(��K����@�{w��>
ǸN�rX�Rzws�{�l̩�3�|K�.�X�Lg;���T���tt�奫��U��5��s�C�� )�φ�=��D2^���
?�.�����96ǳ�^<��.�I��F���8T�Z��E�a���޳_ݒ��D�ʲ�f��
�qV
}��e�씗������s&Tׅi����nװP��%�m�9��²����~ٷw�����8���A�w񪋷��&ʱ�%	�dFX��M�R�u�т�k�Zw��:Y�`�R��I����G����q%�7�.��ķ	��
5�"������c�.��No��\=y/_�y|���<�@�A�-�6,\�5���4�ľX�B����C�^l|��t�)?��:"Z�.�gB�]s;���!���Q�	�IY2������8����'�<b]���X1������>F/��j^����� {q��m�7�*�¶������J�l�n���ͻ�Ǩ6����F�(v�O�R�����`�E����!q�ܤ�6��� 1�������_���W:�|m�Qn�<wFU5�e%F0ӣ�SC��gY��h�[4V܉Cb�_�d+#�^%.��j�t��>y��A>��(�B��EL0���f�6Kd�Q��p��_pC�f%�c'u�D��u=�B��7�����V�>��ڽ�d�*�u�.2��XC�2I���m�� �� ��/,f���`����
�O��
u`#�v��2���#�s+��~�q�z$��r�]j3��j�}؂O�~�{>\�������J�W8aN��Kl[zؼ�Ź����k���C�\\(���:��\qm5��S�u����p+_�U;�$�z5t�g^޺���98�V9"��RK�����~��c�c&��Z �7�7(n&jB�'��w�H�O��ghn[~
NA�lޫ}E�����P%&�c�M��1�D�),|�<�P秾x��,���L�E�a#~5�62�f,	�
���ւ�B�S�f�&����a*[���b4V�r
[��J��]M��(] �g�w�% d��]H���F�8�@��q(s�J>*�ـ>�\��͘�Ae.��ݓ�>�x�W0-��1�&5�X�̀��"I����Ց�W�����<�/j��Bh�A��v?�n�`z��ٽ����k�{�������vk�}�
��������1���-7[��O���E8a�� x�;�ù�Я�EcP�q���E��P��7�r�+��OvW}�����=�6	1�T��R �7rF���1�[/�$��qH�|��7.� z�J��4s-/!%���RVSF�3[φL'u����Y�����&�#�5��/D��G.Ҁ�%j߀hW|b��N=�v�+p:��>D7��](p�ܺl"Y�;��@oF�q� ��F�~���� �uL F��xwa�������T����G�5e�.�����j,���Ӕ������6��l�j�9>��7�i�3�i4`GԷQސ���*}����-����ak�U���j���Oܼ/{���-e�kbf~���'�K�����X&1�9=z�9�yn4��!n��,�I֎��܄��܏�������ԏх�ڍ��:��=.��`:���(.�'�!��6�2?M�\䱾�~3��F���`�L�D��t���������8$��T�H1��1���\�?�8��H�	_s�)^�|���E|LL��IE���۶�!�~���37<Mr�v��y1~��h�g�X���v�9�g��p��P;�}*�"Q;��&���ݤr����q��F�/�jvء#�8�l�����;�QR5��W�h{����P�	�%EtG����ׂ�"G'ň��
�#A��9OR�)Y��"���KcFD�5#�d F3�k��/#-b��=�)�f�)ԕ_clT²֍�˨#4z�j�sb!�w�R��!�P0GEL�� ��e���N|�3Jf�:$!�g��K��7��l��2�	u��1� R�î�V,�Ա,m�A���_��
iQ�1Ւ�.��{�5�֒, #M��	�,b���kK�_3�%����VR���+�ߓ�UTe��Þ!��`��YVè�F���%o�Go�%E �����]�8E�Ω��{��m~�o��=�hY���mU6U�����Խ�Z��8V����*�� ���[��و�,\Ւ)���Wp�����b�HG&��2J��&=���B��P	A�Ot��bY�w��M�|+�s��!��-�#���~��{9��3ǳ�����2��ղ6�E�-��r�d����s�֓�������J>k"3]�mș�C��w�f"gB��@Y+�n��� GP�
7�I̛�n��{���د��y�Ϣ;�u*�ry�Qw0(��;�8���h;n3ru�&~��m�7-k�F���k�D+�`���n�F�d�� ٥*�}�m;�9~�n�� �몊�<����R�-<�T%L!/���Z3��)>��MC4cx�.#�I�����v"7��-�w�U���L�kni䉕8\��ٻm�N���~8'��l��LL��O����I��w�_�.͠Ҟ��R(ʆ >��g�n�RI+��[	�A@�������Ӽ�W�VT��b	��ou�B���Χ| �� $�6�!?�2�s����$�~Gj�u�[Q���C���:3�ۘ���V�a�a��i%�<_��[�l
���l//I�ߥ�N=5
�۸��u��@{�լt��yw�H*������I���K{�S��Z֙��v�K��5li���A�����i)�k�J�:G����"P�:_�N�tc���z�O�6�Z�?�)9B�%��6()*�p��Pe�N�[J�?�g
�	�lS>�#>󙾹��B�A�~�;d%�2�u���t�����l����s���E�}���k���17~�	�b�;8VwR����3��
ǔН��S��:!�Y��t_�bP����.�sϘ�a��%�zW8���3$����v.���	�cj�W�O2���@N�^FL��9%�YkRO����Ra���|������W�V\�1���*�rR��Mc�x�CI��$t�DAE�e��ƾ��ԭ:^\���]2O�k�Ϲ��6����x@_�9��$DZ�o�,��>|U�2˼�+��ӡ��웸��G.����O�R'�P_�����r����Ϳ�����N�{�Еu�z߿���6����{��#MB��#�\Z���l	a��(�h��N��M>��Ƃ�eu�p�f���Ǆ���$��'��z��Ϝ\r�v�9]�[�dL��f���#�V�o~-w�2���G���¨�Q �D� 54�dԆk���w�^G z(Z���`��Y[D�}M�e�ٹ�����O͞��H��)�*BoΩ�K����`MI�W�#�A�e����0&�
�gw�C���1����b��b�E���#O_��~q��Lc��5Eo�ә��^LX��u3��s)��RL2�bOJ�s�F������.\��5;Dv�'&�+�U�1���M9tW������ ��U�^Y�v>�3%��Z��9��O�/�C���tsQ��XX���(���B��`]�Oøa�p�:���:D����j�7���O�����M�q�^�bV��׽�|�!()�<���]�$��X��(v�ׁ4����l8���� w���Ws-NC��/�um�og����Y�g�0�ޣ��'LA4Sq��, �FD���
{��6��������eb��J�z�����[��}���i�� ҫ�Y6�Kd޴��K�ܪ&d���Ɵ��.?���,6B/j �)��L ���-[�$�-�&0��b7sL��У�?K���q�.�ۇ�4OD'^ �r� =5[�쨼 �đ����_:�<���T�x�I<x��BguB;�/q��rK����GB{�f\�?~�b�-^��LǴ29�>�ޖC�/�y�j�k|�M�M�#�	�9�!��{�/@����g��Mʠh	�Y8�b�O�I���Ҳ�n�����J�s\_��'̴���)�p�±n���*��x����=����I띄o��f�Քt��^,A;j�������'�'�>L��`k�b��͍Xi����̺�蠠A5,Y�Fz� ��e��6^�H�#D}ϵ����ƥ7udf!�;�����Zb�����	�?�^2CJ^�vWs����l�AR��| :�tY�0.E�e�f6:1��!��ReF]@�c�,�6x�ݭ�E�`�P�)��a�G�E�I���=k�a1���
�N�)����Q�}��^�g5�*h�NU��9� �r%5䓿n��S�/-�����v���D:�p%�r�����D��$i�����&��
8 �����CA��t�+	D҈���5���L��Y6��ta����D��^T��A���X���?�z��yhZʦ�x���6�8��5�Tվ�B�g���`���`'����i$��E�>��nCY�`��A�\�������=O`S���˝;����]A=g"9dQ��<�C1�ٯX���K�#xYE��g�jy�7t5徖=������J�1V/�1� D;v��-﯏�C��5�E�YcWݟ0�9��Fu���d�Ž��ar�j�o4������:�鬛=�	w��x��q��測���8����p��'\ە���˰��#��{�C�Q����5U�1.���X���X�D'@i|:99��������m뻇��=)��l�Ko	��?#�OW�p�
&��Q�
��P�v˫(�H���{�O�?)���[n[�M�>}�Jм8s˟�������K����������/1��S���(4h�u��r�t��Hf>ϔ����y]Rn~t�žk�n�*"����21m�f��"A���b6�Oc�hK��5Ő8A�F�JMշ��6T��3��|�^E#V<d.�7�\33����M	K��!�X��ˬ�
Y�æ�L���$�^K���Io1�ۮb��m��(V>�|��L�������=���M#��Ý�e�F,�^�p?�?֓R��v�z�=���(UQ	�5����*[��$ݺ)`,h�)�BO�J>s2	=m�%���z�Yy��|݊]�D�rhr$M"��}bct|�F�(l���1l�$�����\U��}�A�vW�*io]"\�9v	�Eo6�d
�����4��?2��_�~8C���5!4����{,�� wI�Cִ�o?�V�X/�{���y���q�����5X��7en�dF4(�i	�ץ�]� f�J�teEkh�l��T�$���i�|r�Z`�y�T�$�iI8�H2�_t4e[��&	�ך�n�y{�[��-���tv�`ю	||W�&!i���$#pIn�
7�/9���c�	{��R�Hin�(%b��?Ɖ��>q��tu-�d���p�-�^�Q���̓K�25�uS\���?=�`�3�4W��^�"�Ax��x��-��Vph�߷�����Q^����K��=�(�=�V���IlYG��Y%�YX�
�O��:	E�j�}$
�V�˂R}�Bcjz�^���SJ29�v�ϳ�c?6�}o��yET<ϝ s����4����[��ڹ��L(��\�\}��-Jt[��.L�=5r?Ӎ��}=��@�����?y��Jbu�!�W%9��o0t�ڷ̵���l���[�����~y��+Ig��H��Z���ƹ*5N0��jI�.,K�0�rV�K;�ke������-�s����H��&EJA��T��3D�@�����E'���P�Q�S��4��L��#���%�����|����E}w�rҫ����b�iw��4ߊ�oFe��L�bL��[N����	&������4o�K~7�]��*�y�������).⑄���h�þ:�#
� zA[;1]�݋�����`�[a���rl��'���c�
F��p�$^�k<**q3G��{5�֙AJ#^�D�Y��E~y��q1�'b5�b5�<9$�������osd�m���4u&O/o��1�=*^��+�}x~~�^���]�?b?�vЖ��W�^yI߻4t��Tǜ.�gƾ��!�F�JE}h�|/p���R�����ʏ��g��si�p�V�|�Ʈ��x�J�����"��g���y:�)�f�Ϣ
�H壷�E�]�� ������
 �0?�fǠ˱���1N/�=�Ase�Ϋ�%�W���W+�;Y!��w�RE��\g6/�*^��0��[�����Ds��	{8�vY�Ù�*v�zL ���8^��u�Ȑ��۟����@�W׻,H�/_+p_.����v�,>q�tc���Gዣ#���M���&�ļ�6��[��s�po�+1"�/.M�n�z� ޸|9�R1 L	+	B�x_�3�#<||"�"�'��1 !6�����+�RWL�bMx~*�66d�~w�hb��*�4k�	Ʈq�h�;� k���������@̗/)�v,6��'@��L���]�u�n��By�&���^�OO����Y�����X��!��ExI�N���>k�Qp�1.���f�3���I��Oko}����o�Ktt����z�6�J�Zt{��.Z-���'�O�d�X�U�}hx�0�X�[b8�/ �bvЬ�J/�v� X���$a'D\�^R��,8�_"�5T3[h�?��W.�q4�)8.�J�n6���Nd�=^�R�Vh�RǇ�ϖꜷ^ƶ䞽|A�aF�	I�d�&�Ĳ���18p���E5��B�����w�~��`�^ �?�s�BCCs�N� �)�atd3@������U�I�e~b�5صw\�0̡H��C�J/:���(_-�Q�%A^CJ!I�K����S��.1	k��Ʈ�x���[
0��7B�j��<��ᏈQi~��!IIM��7@'�ji���<�������Z�4�E�>�|�L��[�Y�ǘu��z��bp�E�<I)Mc����"� 1��3
		I��В^��~NT�+a`�c�>������. f-�,��Xh�,���|�Y�v�^�D��9`@	�=JD?���_�W���1��&��Hi�
�
�k�Op]��F�T뿣
5�EH����4>�t��φ�S��W����(��Dc\%r�)��h�w?ܹ���1M��V#�f)+ h%�_=������T ��I```�����)�x�ŵ�O	{W�!�����,?�����[�V�#�|=�w�;�2�'
��̍�Z��5H���H�� J368r^�dQ[-��� �����鿲b�oj��)T� ��*�XKsը�w(Q��8y��`SB�+��N@���q��vX��`�g�錮 ;Jӆ�j��Xc\}�IE� ��$m~�c,hh��� ��@��`PX	 D����V��c\��{���/g�胢��O��
�sČ?O!?������,E�ϋ�y�C(9B>��%}`dDs����ai�\N��}L�����	a����c�>�b p��g�xΰ+#c�y�b"����..��|���<ؖ5�id2fu|m��!�6��^g�b�[�B*J�ZO���Y#4�~1��&2q�+�`S<�g[��z�яB���r�C�~�T�l�ʉ�B�b7��:� B�s�������	�#n|�J���x���y1:�Al�b��g���&��H;�D�������
CD˫2�W�8�J�����0�h�^��}�z��x����u#Ϗ 
��l�]�B̳�U=V	�cO��J�9_WY��P�/�`����J�
����R��e���;��yFP��A�S���D�ճ�TU�[�����F7�8��=��<]uXT����F��Q�^Z�n�{��FiX$E�;�$�AX�s�wW��w����.��9��9�ܙM�~�!��c�!�Kt�x�(��\NV�o?���p��r�'�Y��l񰻣�J�u_�M�lRQr�7	C����d��Q��#��{9o��4���k�S�9������F�B��K�0o��Ð6������1��49-��Cȴ�9G��'%�/�@Ex���pCe�/*�.z���2���)1�j�v��+8��� �Q���a>�q@�@�YƉ0n��s7��R0�Q��t��d������_��IJ0�D��0�`�Lr�������z���.�2���RiG������Wa�H\�!WEZ�������c�=�EZ?�0ς�s\? �_�Jo���H�]RJ��v���]�pYy9>���۟v��c�":��8��ۓ���;Huw��o  8���"~n�zP1;.G2"�rʆ�4�I��W1���@�+`B�Y!�c�o|0��(�\mE���5cl�910���p'/|ӀU�,j�l�w���R|<]�������L�ae<�#F�P��:1�-�$ɶ2���Ʒ0<��"��G�_���&x��V�A��b	ݸU�Z�#�~������=?0p *EXd#0K�X��2�O���s��Miٛv�T�}�T5���1m�<9ۈ�U<�>p�������XU�Ԛ/,��#OL������(��C�>�񺟾:��~��J� �42�1�����TV6�5�|�z��	�<$�����d6=�F��0��$���BEX���:,�KS������?����_��-��}}��|�vI����a�6���!|����ge(��`��+ܦ+Ъ"T���w�w`:�ڛ�v�p9����µ%�:qJ�+j�ӛ��BL���� ރJ�đ���zx���sT{DC��8��E+�Z�D`hEzq�f5���.����) �X/	��{���-��N�|.qy}t�	�5�ZHx�C��a��_���?�ҿF��{�,�P~��è$����B�����I�aBV�=�V��P����{C|W6�iK�l����ơ������a��w�r�p�%U�997�=�tf�_�b�e�m�#�A���#�w���'PF�Rac'��ϊ�@�%?�2���˓܇�ԣ�h�B�X��R���ϳp~6�W�&o���+Am2��񂣚�~�����;J�m�Nl��~�[(adZ~���V?�h�ewa�d�-�dƞC͍Ӗ_���(ϙ��SÝx4� ��������^Ի�o@r����
���zL-�˭�"��3����}����\��s�}^�]��:��o�����/�:ӡn	�˘AY�|kEe��ɱ�^��������mE�N�"�Y�q��K��!7D$Y	���0��MCk9t��u�>���|c��E��#����]�-�&�x�>d�=���&���wH(�t
6+u��iO�)C5R9�H6Ltw�����UJIgIY����mLcͷ��\Q�e�	�,�;Xr0�GJ����h�Hwcw���;;���'s>��[��(�&P��@h!J8C������g��j�~�բ��6�Ym�ve1�lE���D~y���>��6��g��0��6��7,�Q��,@����
�Wb��"�<�3����~^��n�0ʽD�1f/�ɰ�9dw��hݯ��_�(�܊�X�M�[��[,ZD�|���c�X�2}n�`/ALAII	�S�ݢ��V��$pP�1!.�����Nxx-��/Wh~��௄�|�L?<�׼��]�kp�J/>�J����Z��ᓕ`��R��-Rr.�rr�!?J!&�r�J����P�q>�6�������p-��~{�we�d<�婃��(��*��ͳo'Ȇl��d��Mk�@>�9�3 ~x�8j�=}�8�����N"���XB�q�]�� ��{9�q#��sfX�}���"�R��I��$[�Qem�����v9����0t&��[�꟏T��ʾ����<6���z����Qp'���ѺAQ�8�X�jY���-5�em��R�js3N�S��O�NN��iD�?I�"��bm�<�}�a��2���,�*V���Α��U!�0�ԟ}`��R�ۮ��݅�2���0F*�D���6�*>Q;Ê8�1�s�*��Q���ܫ�%^�_L*5Yypj��x�;̕��-F����r�����e�3\�s��Z%K"}�jn3�O��z�x�:���L��h�/>�Z��z���0-!66v�u/���=	�h�.���G0���F�D�ø�=�R�>����چ���K{"_ݵ�*3��1�s��˦0��˙/�fT=�7��~i���"��ۅ1��ǎ�TM�h�3���}�;m�r)t�"0�\e�3�A\'�"[N�s���[ �S\D{�B���o}�D���6l�V?�!�E���ܘ�Nዉ�8z�k�Qn���D^Ɲ_�ǁY�3d�@�� �4i@�����gZ:�~¯��K~1�M,��Z�>��[�s&s���İLb�Cu���mƓ)�)D�9c";�==;C�ñ�J,�����a�E��7�C"}�?t��4� �+΅���Z==��Jy'}���Eqԁ�gƒœ��I�v�ȳ慿�����s%����~N;jcАqϞW�4�ȋ�j9������8�ZN��aͻ&D�=aʕ�L���.@�0� TAm��D�o����0Go��;�I��z�Q���)��!kC��:�j��
�8�L�r|_p�������׵����<��q����R��p��9Ҵ�b��ȤNA%`F�J����%���iqn����\�	#ɓ�1:�>�.D�]w%	����RNAD	3�r�Ԫb�1���!�_V�%3��=�iRw�^w�b�g�/(�A�ֳ0���v2�b���5�O&=�m:����D����HcD������a�}ּ�*w� �A�4�����ȎZ�T�`�P������II��H
v�_�"W�S��W=rO<V�Ը��L�{q�G~��ri�%�l�)�"�,b��~N��
^'�$���.��������#��<X�HJ����%\�"-W��#M8��7N#�!O&�M�ր�#�թu
;�Q~�Ԋ�Њ��+'��DR�u���h�Wq�~�X�o�n1���x:�'�|�,.PB����i1��υ>z�N�y����z������LW/���~�Zp�0��������[�&�kZq��M��x6H.rUG�����RL[�g�-८��H������>��GF�E���E��S"���晑���g+>�Y��6�ղ��lj%���J6р��m4h���[`�V�X��_qhk�\���`61���Վܰ����C��Ȓ	�?��5�x��5��b�:%�}�#H%��V�5�{�7�cH��Gb���7oWK�_���j2��pR?ϰ�'𢣬T0Euo%��������<����M"������2}��:�b?[��E1��ت�9T(��Cr�^o��8�:�]ot9�����A@���tY���(�wj-�;}B���^DU����������:�=��u���  '}�_��	2���<].D��+�Q� �����=;n�8��1�|�bR�^Dr�4���ˇQ˛Qˇa���=�Q93�c�W׋�A��pOգ�y�Yyuޣ�O|�ӹ̩�z�s� �ޔ4��s�#��
�oi�s�(ZB"*4�ԩ���G�qۣ���yA*���dF6��7��bȋ�u�d�^I�I��Lϑ�hJ��kL��^�W�1�n�n�=&9��,�P�V`��q�$3�vJ2�Q�"&Sf(|���k�)��4���r4�o�����:Ar�bK���  7pm9��u���U��_��)8z;!w��q�W�gp��>56OMQ���%���n��hq�8�pG�<��zW]���HM�T?k4�"+����G�����ͩm�PD[��i�4܎���Ta��;�{r�R���}|t��#:q�u�I�������1�R���	c��{��Եx>�z@�!r���R���5V�o>H�4�������f5�]��ZaUL%2_����!��:����'��Vq�8GC�k8)�������RUnr���)��2�F��N�4������?��D�e"����~�8���t6����ZW��*��	�T𜜈��F'Qj�/��-ۚ�#!� ��l���6G����R�a�eAn��=uS���+�H�� �2y6����Z�g�M�d�� K<��/��n3�� 
laNoo��Y�����ul��0tLZ�+B��혏�n�!J4��QI�q��x���=��)�?E`�c�0s�ӹ�UIf��}'vSq?��~�ĝ�WW��.X��ƾ�|�~�$���L�ɲa�t�(j芀O��:�&bǜ���_*���})p,��t�Z�՜z���_C���<�vx�X@�ĉ��'�Sb�kaa����C��čo�Uq[t���+�g>��Y7؉Q��ZJ�˵b+��1׌[�/"@�G~t.�_N���^���E'j�VT�
�pwx�B���E�b�^���͏���y��DJM9���CJ���`;��:�T�x�d�]x��jY6���`��J�1G^���8rO3$`v� ?�7l��3�7A~�!����;�<q���C9+6~qD�9�ڢDcl3�q.���-� 0�c��Y�C����+:��y��G&UXt,���z�#���ɠ�����ubCO�#���6�q���ZF�c�,�Zjua9�V��h������e��t^��(s������ ��n����d�[9��?a�G�ѭ�<V%�w�ί��}3L�V����`JǾ;����OF@�!H�TJ�A���C�Kf�>���x��pX�=��M�$0�1�[N�F8�ѓ��N�w��-�����c�����z�t8Zx+��9-~n`�G�>5�T8G' j��t�-X���	���3:c�IΩ��;.�8l���N��O.�T�p�ϡ���Tt�1W���p�>��s����t�� ����׭wX�����|�o�H��s(�⻊����Q����K|��[q'V��n�$G%�J1��7���U[6��&�σ~L��
O�*tj0�n���P�\��m@� 
���'y���;�Ċ0t��ix��q��}����Y���3���<�k�����e*fG<l�z|.b��R�`Y�ƃ���Ʃ`��l�{f��su�n4��u�����lϊ���{=�dm��դ�� 8������zE�N�_�Q�"F%�q��^ɾ7?��S��c�a�a�P�L�aj�2�H�"剌��|��h���}羣?��!w�b�y����i�I����PT�AA�i�]l������1ee��0M���Gs� W�e���ã���1�~g�R���5�e�8��G����=�P�1������Bk�%@���v�(��4t5tS8W��C{�A�c����K��|�rD�.MD~ ��hS������~Ӣ|-�3��!L��I�ˎL�R�@;���s�Wd-$w2&QUN����S� �����j�ɸ%�{�/�q]n��H�u˶�̠�:&�j�z,���D�/~��.5�g8l^�Q�:jjN��8�G��Y��~cT� �\�hՖk���ۿZ��
v8-T'����R-}u(�;�G��d���3�7�C8�L������cu��x+�e��u�\ő��-�x�+q�;�
<
=�w���ot8X�{~(�I�J��ԩ_E@ә<���M��������tC��e�^Â���~�I_���|��d�,�;β�6�AG�5�b�j�A����Y�є���Vk��cU�p	�d���?(����C<�$r2����ã�]eׄK����-� `9�<364CMCA�L0ܒ���I����Qq�����*N>$v/����J%��f��=��M.���R c3j��ɐ��kڀ��7�]��?�7�xq,�p�B�G��BV6qi��j�$~����%@����r��|A(�iD̀XY���ލ�)l,D�E���H�hr=�_
���p��M�n�ݞ�$�����q4.Q��13D-�7膄1��T7k��*	�~,#�f��z"δ*����.���w�#�=fJX�Z�<�����6��f��E?�_=�����˙�\���[�!ܿ�X��9�q�zI8Y�px��ʉyKK+E7\�	T��Sq�O~�)l.D�U�6Ө��Q5�����El'Sd��wo���-ى敥�5K���{��ZB�q9�.Kn��mΗ�db��&��C�6.U���)SD� �����Z��FG�-����WP߂�6��R�G�Sv���F�(.�G&����[E�3S���0��0��L%�*�
/O7��Y9�US	���4��yl�F����2kx��} 'w�����	^\�ITO�S��$�^nr������{�ـk�O��ē.��*��xu)��`c�{@ǇW�!mjZ%�v�8ŭĚ�h#BsG��K-���k���
  m��:�E����}b�!��u䟠�̇U�4�S�GW���x"&����r=�ߦ.X��w�C����/�����c��e��O�[xm�Q�(�ZNz��r�R��j�<*k���u��O�"k8�Q?.B3/n��Y��[�Ë|R~�3:G�[M���5�*�<��f_�¼v�Cr�����N3��u���=�P���g3rQ�x�T�ʈ�|��� ��*D��6|�d���j!� 0�[pcƠ�)A��|�i�\���i�׸�Ks�3'��{���P���x5i��7��b5D��s,σa�MbD�l�Z�zT��+�/a�o�3��'��S��tָa2��_	S�RX�4��&��)�IE߻�}B�L�Z�e�^�#pł�Z���8�.~������Ս�Ip�SԿq�|�X�[M��������R�����NV9?�C�{8(�&�6�� `����¤��-x����`���6x��щd����ӭ9͝?�D�!����Ų�)�=�Q�P��RY�cD�pyD�5{L�0�G���e�p�$ż�#WR!��b̏�m�Kxp�E`c��A=o*����L���ǈ�����v�x�Qb��?��Z��`�Pg������yo��Y+wE&�O_�uG�;zb��OI�����T��eL�ȓ)C����`���7�JU�U�NH�߫�<G���nU����r��W�<�$W���	�,��X2�M|īm۶%ԃv����܉����`���'��H��MJ����ᦈ_���j%�~uw�.��ƶB��7�Ż-9��%�����'3��{��8��5UJ|x�����cO�!��x=��H|Ч�IbG��j��TF(��Q����Lt�+�bԊhi��e�esū�1�&D�"�kX|���[�>��X�\��F�W��p>�#�/��.1�q�;a�{���Yӫ��ɤ�ݢ���<�8�\}��䧸�R��4|�TJoӖ��d#O��t�H�f�y��l]��
��k���ebf�C wY��7�1�*mH�'3*�K��l[�k�+9�� F�2����K��*�����,n�X޽���fB�N�WaX�=KƎ&��#�v�O��E�mrDˑ��YrDD�y�;�+���2~�\}�V��g�`���%Q�=��)�߈6�N�A�����3 ���[b���v�z�ʇ�$ү�����lL���ݵ���&1`zk�n������4i%E���lf:#�i��k���{#�`"��O��d�CR7"�6���C�>u̇5�>�3�Y��	m-eE�xJ*�%u#��ߗڐM�u>wZUQ|���v�J�w?�L�ӱ��F��SO�e���^�l��ݲ/�=w��z	Y�?�jS���K~�`���Ѭ���*�wAިo~�,#�� $=��}��Q���KA�O<�bع~w^x^{�	T��9��Ű�36CRlJh{��;T?�ʲ~�ܴ��.v�����!�r~0*��ߕ[��
��Ҩ�m
H��`�pW.�w2I�d]'�p�CG4Cno�kJБҌɃ°�d��ę>��K�۝�ȫ�s�j��+IoW�ؕ����S��-�+�&�(�A���5�j�=�;Ҫ���v���es�ʯ�RU1�q.4S��vV
��aM�e�	��K_m8�UF�9�(�i��gQ�TX�5hsl�)���ũ��.@m��f���1n��b{j��r�&���M�QjM�LU�g4ϥ�S�a~���j�J���]>��%�©��ī{��R�|��z�ę���W?8��W/Z�ڊ1�
��|��E���}��i��>5��4�~)��o���Locrr�/��URk7�O����(�Z��Ԝ�b,�/ȕ�}r���f��T;wSl�v3f��]oY�~
w�����0��^$-v����,ō���@[ɠQU��q�)S�����R:lv�\٧t���מ�G�
���<o����ҋ�4�/�R�#Q�ʖ�g�n<_�b9���4�713!�	���+\S���l��5�0���Uu����cI�D~~iI���1�|��o�K�o�j?�gr>lZ6�Lx��$ ��4�lk�0��{�_ &���|u6����>�qOZ1
�7����&)���� �vva[<�_ʾ�UQE?v�'w\�Լ��v$�z
�E��^hu�!�'�.�[����5ݣvs�^+'��ç��W�e�֡���M�jZ)��\:�8�0��z&*J��H!�&�D�L?���L�2?�8y1�4ՑWw��K�ˊ/4��������Xni�h�B��,6�4�΅�B�a��eHgJP��"�~�|���K
�W[�X�Ǳ��}i�w��\�����
���)TO�,��>?��M�ux_���9{/ޟqa�9W��r��T�7�Y�>�W~2K$.Q?��Y�!���x<}:�I���a��>ALU� Fh�=������
� ��=@�l-cԍ�=���0)7���>r��ЩW_M���!s��zG���]�$�8BĘ��4u�4��(�[�9�U��� ib�|��O�����Xw5���]�D�9��Wff��7��	�� �����fu�o�dT�7���V7Iճ۸���X���֚?g�c�w��Zu;�
r�9���Qm�-$ݹ�nD�]�ϵ��+}ɠ�� "�$�,�|�#
[��]��f�Cj ��Ja.���V��6Kp��	n�����2~%@L����c���������:�,�p�Sݘ~��pxhfp����{�k��Q�nq�Al0x�V^�q�Ⱥ�����O����H�x��מ�i��m���w"����s�K��G{��C.�Y���!�5/dN�[������W�~��H��覾�f.��g��t���TOd�L������	\��y0Y�е�A�)��op#���y�}۝�q��?�=ҋ���<|m�\^�*��q���m=�j���QS^l����;�pL!�� {+M��գ	��4'�I���#��b����U��i�mȃ2�K�O��#:��Čvқ��s�����.�wЏUA'`��������K-ߒfx���xV�����p���~��t��wBȠ�������;sm�׷��SFyʩL��DQ��H��?�{:�:�w4<����'O,j�_6�����J���,5]ܟ��Ӹ>��A���n׎�/�ʹT�l�aIha���y��UI�m�R���;u����+lՄ����|�v���uv{۹���a0��[�M�.�~�F)y9N�kT'M���e�>U1$��(����7{u��s��gu籤�^9W����a� �N�Ѣ�A��"Z��I>�[�<;���S��,�ުP�p\c���lZ:`�F9`<�������y��0 �;�rf5�O@�cJ[VD��U{';�w�G��[��#����=hd���lg>I�l���Y
�(��W*����5C�cMO�g\j�!SzO��*�^"�#�aГO��t3����9��K����_��Z�]&`��Kv���1���7��܆b���:��u��\&�~±<�����l��U$�����n˵��Ec�����	�H(��J��܌c�˞�1���7��Igs;e����/�N��H����H������S�m{� �U"In?��nd�@�23���5���4a�{��P`c���[ۑ*����$[-ۮ�u�%��D�>�x�#Iv��K<>ݕ6R2��v'�m6%ܝ�e��C d:��[�3���/���lo�W��(�#����5�b,��ߖ�]V�i*��rt��Y{��غ�r�G��lʉ�4^�h�����������3�hTگL1�ع:�K�UA┋t�ڦ���j�TZu
>h������K0c��*2�;~�W�q-��$����-��4���甩Y��O��E�@J���i,�	 BB.�K�Y6�~n̳�~r��3Ӥ�@�Cr���Z��7Y54wR~�Lh�E�/OZAB��+��-���`�M+,AWCBw�����׊��Vm�ҜX:��D	cL�)e�3�<�^�.���kQ��-���Sێ}%��eh�p^ʯ�ݚ��}8ᅶ?��o�y]���u�q3���� �������E����j�0�L��u�ȁN-`TYNrTHYC�%3|zP	�~��IM�񄡞��
G�W��/�ͤ�D��6�D��+�B@">�tޙ���#��4;�P]�~u���~y���	��E�q�)O��n�;��߭�PX�!��>4�ϗ�Y�P�4/��k��I�!�^��o�bO�B�1�v 7�'��%[U�����7ꔢ����9��C�o�/�'�;�"�8��jU ;�eն�b�����*
mN�<�lTL���5wm� �@~+�^L�D]i� �N�=�H�$2Tt���O��G����,�*7��sTn�}۫`����,&��:�ej{�ݹ$��o�T4��&c-��79x�oq1�mA��Ns6zC��"�Ê�bv�������kM3B�\k��A�ϱ�*�G��&8V:s��3��r�rf �O�.��l"Cy�J��8oM��t���}y6Y�7��+n��D@����z/�{�?�D/�7��_=h����v�iЅ��!u�Wn�]վ��A�
���đ�0a��4"��g�9���jq�����"�٬#�>��]R�o2�<�>�@���m�gn������ŝK?���	Q��UC�������䝷���;%����Pnp��&����(nlF��l�eYhi�-ڵqOTNu�2�R�S��b~�Fb_�M�H�/�6�m��������8W�a�Y
CdoϿ���\�h^x��r�5��3�ը*3�E˛����KR�Qy��u��L0�17վ��
���OW�ko&����?�0ÀT��_T@(��~��7��i:�8._:��`����;}�H�o��)���'�(�gz��LEOڨ��`9�pǵ3/��\����[c�㱊�|_r�.�u,|e1�M%�68ј�[~�!�cS�gj ���:��?�$�O�Z&��v7�b0n���_h���B���U�p���j�m�?4Z�IY5/��R��jIF��ED�Ugϭ�~�[p�̵���@-�.�ӱ�aE�;^��m-A��ᇉǀ7�Cy���~I ��x!�%N9A<J�GR�?�
������]��������Fbc��W6�9n����}��u����|5aH$BIC�1��(S0�U6�יǪ-�V2���g��bf8`|h�����J�����P�g�3C*w� ��7���"�һ.������tD�R�i�'nB�H���Pm��X ޱG�L�C{m7��qE�^q�x����y�{f2}|r/b���?R~�/�9�O1g��AM�/����H�q���4~�BN�v���}]�0{�`vJ�%Ƶ���	fzO�Z��k���j@����
n�y���vu�	��LM�a��g?��KD��e��7*�bI㬠����II�$�L1۷&|��C�%:cx~"���	�#�8a��L��# V�	��4��g=n�6n�fǰ0�߯ܵ��\I�-��B�y�	B־�L����vi%'g){7vB���]��F��O��<FqCD{`4��}��Bͱ���2�l����tF�s��o���ޛtj#��nL&�O�^� M�V|#��� ����@�.�j15,��)L�	�]��\;�+���G�l>��E�Ok���� ����	Y����2�\KR-��[��)k�G�2����w07�,c!5o�����Rʨ�D�������(�f�.�}5l��8gp���c��\`S����*m��x2��my3��������&�h#���6���[y�DB�Y�UQ�A,��0[�7�ׯ�\�Bړ;�&yQ�0^	�x�� (;�<�3T��VS9\z�0�U��p�ҷZ X�u� ��r\��qg�P�g������<TU��h���v�wWI&��cP-�1yź,����a�(�mC�F>�%- (gn]:ea�8ٱ��!�g���Rߪr����ĩ;��p,���v�������D��~���lI�뤰��EN�e]	�y|nfl�yg�Cr�|<��nk���z~��)7���f\�B�]&z�E
^��׌J$3-w]��'e���[�:j�U�:gKZ�NȐ��o��?0����c$Q��#����u�?X�f,�9ǣ�0�����%����㈼+�u�k'�@<�o�TWt'�XP`m��^�}2��ALe���L] 0�)��֚M]qfu:L�'("՜���IE���M|NX��[k�ᘟ9����q�m*���<,AS�?�SrQ壚+�g����k���M�e/v�*l����̀��:0Չ(nRCmS ѺS;�Oe#��Uh�={b��<.��}�G��&�����e����
�e+ϟ��>==�G�\�q�)�Mr��ٷ
���Ϛ1���]#�Z|	��\J�)O�]��*�S�nWC��؂SUݹ޳y{�G.ϲ��?��"�7���u1g��z^'E{P�J�뙽�7�Y磥;m��M^_g/����ߚ���i�B�B�#>Z]e�Jqҫ�w$�q�ZIi"��N�eB�I47���-�;y`	��r��C�ŵ VU�y�F�dJ�����5Y����|�ɼ���>�~52�:�E�7�Rsaj�ɧȪ2 f栖]�Ȟ��qn�=A�-��g��o��D��<���4��_�.�w��3�����D|����ti6Y���C����ŴҰUM̄+�%-�Hh�@<f=�k�2�2�Ae�`H�9�)Ѥ�E���T��ٷ9JX�l4sA$�G��Mkz��V"�y�ö�Xl����GҶ� ��֛��d���d��J�cW����7�@�[�"VkP�,1��u�y����;���Gշ�Z��.K"��J�f6���H�1�ȶ�#��}5�(�"���s<�ޞ�d�O���Mv�~��җ��{�������/���f��`"<���9W�2�7��o��7��X̍�|z0���d�?5]6�#y+|�T`�01Zh�8V�}%�ͳ{�i��	�Hr3�n}T-���Kg�:�wB��(2�Aԃ737�M�*�)�^#]�3 `�Q��`8��=�i�)x����}��^lק���O��	�\����?ߍ^�BA�,����:���֬�V/^H�'mZN�u5<k�&�
��39��G�T23�E]a�i�~s�����$zOjӒ�W4+�/��P���ڃ�Ya��˔�OL�D��{0��$���X�טFͲ�~���܎�p�\^�S���q� �|���jVƆ(ٖwCeXݥyK�*w��z�kcP�?)�zDj�z��`}�ɜ�pk�c�$���f-��a�h�"��H��N�=��|v�ZR,�ܶ�)���dlGJo%���m���/�)S���n2�2���d<%��q���D��EF�����Ǘ���,�B�a���Ǯ�ټ��f2~1�f4gc=Q���s��xd��"�i�=#-��ϫq	����{X`|�^`�-/5��%adE�������ۄ2�i�}�Z�$N�ۘ����x�E_`dSN�������[����;�D�T��ӵ�l�R��P?��=d�eJM9v(ô�W����_}K��T�?Wf�_̬�ޭ���*f�w?Ҳ\&���Ш��Ә��=��L���=���c;��8<MԠ�S�o�ɶ>j��^O���/�ѧ>�L��a�3z�5���!��{����e��a�T�S�0���g˜t΅ɻ��>��6wF?��PJ�	�JR9͡�$�>XI�+<W���T�<ϭB����)�]�oR�)fƓ?�rYQ�0�e���v��/��Q!"�99��7f�]��<(�\�����|�Ni|~�t�`#�`����{|摓����Qe��{�ڮ���a~B��Oi��V6pVc*�Z�,��E��*#i����<��������84�0]/�M�:���^H3�?3�}3�{�c@+�R�b��ݽ�}�jvDeT~�w���>p� ��2��o<���%����m F{�5���`����j+'?[����qC�u�!t�<j���Q��o{��,�/������m�N O�����̈�� �,�2�;+�C���?跎�~;L����,�L�E���PBeo[�v�o�&TI���U^Ni��O�	 �b&��ٴ~��1�M��)aEsz0b(k����]B�9�c�z�,�Wx�D"]�~g�S�5��g�%4�ᚨIbg?\�1 q��ͦ��7$]�Of�<��{�|��<��aEZF���ί8[�'8����: ��"a��Kϒ�/�G8ju.>��8C�r6�:?V�E=�?v�R�����
:V^�E�=�H~}`?�_J�}�g�}'��_�xT@�ctS�<������Q���@V$$R|��)���<����� ��cQ��R捾ʮ��ߙ_{O)*\E�u�.�=)��D3ؑ^��(�r}���(WnC1��..��B�'�r��"DѕF���+UC�C����@s��+��q%^��<���;�֯��|�>01$��n�;�AS�M��Aţ<DT!ӊ[=�7k�$�R���l"ϊ�a��c��Y���D�[CɄ�vJ�i�Q	�m��&��@9&�?h��W7�={���^$LY�i�=�D�zd�{����(߷��9����Gug\e�v=��R�ν���O�0�(��5-r����:C�<�ޏY��ƺ�փ������d=����.�D�O�w_�i����0_�ɚ���4�����܂f@,P�f�!5?L�}�ՓE<t��r�լ�E���z��� �7��:Kr����1a��z��.�|�%joy.��v�h��ML�U�Y��@�7\�����Ję$�n����������A��^+|��B��_��o'�%�l�}�^�(bң
���:*,'U����?�L��:��b�t>.Q*-�S?@O~b8�6���d����u?j1�Jj�V���U�}5���,�����2����{�Jd�ٞ���"����S��դN�AE�v�D����mR���H���>3�[N���Ӭͮ���XZ��ݗ�y�i=1`�!�ظ2&#��%ip3~���C:�q��w$�IwE�1״R�"�8w��`������m��~?[�ܬ�46�nܾ����p�9����V�qu��U�f�W�oÃ�Y����ՙP��9\�X����S�`o���p�.��GU�9�0Ύo��1�O�Z<��1�~"�l@��j�^	pP&>�b��z� H/���e�Á%�fd~��?=S�,�q����s�G4e^Z�b��BX�vc��ֺ���[Yﺶ��/��1����	�](��,1��m,�N���p
����5�;��+��<v�!�)M��8Ȓ1>�oճ۝1�L�h��ak��&�^5���}���-�q�,T>�I"�n?�)�L�,@���ؗ,r����
��
`�#XQ �H�*&��D'J�}�	��B_�����^L�	�RKؿJ)�$��L�!lt�ݬ�^��+R�%�"=1%����m��\/n�X���[кK$l��N��RS>�!B��RдB�{6��]�۟x�U��]��=�k4W��O�7�nS��H���Uz��UDdvw�@��T�Y�*}�cٵ�����Z��coc~��ad��^���w�\nJy]�yfMm���o� ���'��
T��0�]kU����楅i��r2�]�Y��V�J�#��4z�;\�Yj)�;��Y�=(��^�c1�JOt�2]P#L��=�ظ���:���6��6BH�Q9%��������u����,�p[�<ٝ&�Zr3s��U�m���D�������q���nvM��* l��cͲ(���h����1�;���
��mtz�to���#��u����Z�ޑ�N�>k�*��	����lX�}�W�]�ceC��1wK��UD΢f��=�ܖ(Dg(ߕ���wR�eۚ۳�FX�+�#�J��v�
4#?(����B�i������խ���nd1K��
�n��������7�ի����㘉�Wqչ��Aϳ�_�|%��+�Z���W��Y2�.�go�5\�p�w��7WG�R�99�-;e� /n������Q�{�P1�ը90*'��w����?���-����ni$�KJ@�AB:��a�ni�eH������!�j�����}�;�3�:���k���9"�3�m�:&�wxxͻ]����s�b�xBX�pF�k�"|�b��}�|�g�>�%�΂=�E�'�S��n�ٔ�����]�O��ĳ�HlTPG��w��VP�l@��@��t����tz�	����_�7h�����6��+��Nb�dak�ǝx�&K�v_xJ��:J�.2p,$Ҳ�p�����X_4
|f�1-��������o����C�Ә7�v�;cK�;>�rң���Q	r���@��J��2��n?!P'��*�C7�A0�#%$�A aTY�����VQq�Ft)N,C7�ǲ������%��� ����\-��B�I/�����[CL)C	��y;Ѕ��X.��(�5� �����"�u�AA��v��R�v�A|[T;ٳ�M+{�g�uʒfb��A�vZ\��������X*�7��,2m{��Fr�U�{�Or�0�y0:���Ȟ�S�n+���츎;�����2c�U1&(�*3@�8�G�}�6�^py�f�]u��q��zaOY��h��F���Ʀ�{2�����#l�m�U@�>h?W���@7�À",��y\�g7#�_�ĺ��lB��Ck-¡�OI�k���\�{s�J)�Y5~_�{#)u�Q�\�I�_��G��'��%c���+@ڤ,F��'����*����3��w+�y
��?�"�x��.�{�`җ�}�1Ok���r���װw^�!:�����+��67Y-'UԠ�mz/��p۴�hr�;E�S�v�iz��6����.c�b����cU�~�ɳ��a�M���|��c�ɾz�P9�\P�E/b&�΋Q�V��{�cmF'� ��wy����ۂ��0y
W�m ��M�g����?{�����Gٶ�6 ?�}��eL�z�B�kU&�R��^:�+�d��[x�[8����3����ُ��xx܋g��0Y�yF%��T�0�T��/��Y\������p�F��elv�k*&ç3���'	ϡMBoŗ���z���;ڿ�0^�����NI:�
���5�el�9(o���EgM��F������ݑ�s!k��o�;{�?
ڀ�"��:�ñ�������P�X(GG�
H��}Ds�4�͠M-�F�ҴaD57v^��A��8���� ��L)a��S�H@�����s�㫫(��deޓ_�`)}�7�`�mv>���!ΕU�1����<��7ܳᤶ�B�q�� �)g����"QR-�JE��5��n�R�Ú��������NW3��Á4�����V�^�x�^���lȊ!rxK�<[����%��܉�Ă�������3�F"����k�?�~�q)jZV�P�౩�ݬ�_y)iƆ<.#!�ƀ�_H�����I�_d�
)?9#���������sj4.��t4?�(ͥQ�B��YM� ��i��>Au��h�|wȩ΂J��ɕ�ٿOF��,.t�����盾Rف7o�'8�0��JPD�y���Ap������J|댡T2��:o�m�HSߠ%��}@�Y�l���/����ا������k���i�:Un�9!��ˡ���.�9H���ż�b�o�|}��n�,l�un�)��Mt�8YOU�쀂��!�R�V9��7�w�E
ϔcK�Z��a�Ǘ�e�Z�Z��!�ڧ�t?V��ȫއC��ȅ��{E�z���뺈�wh*Zj�v�����0�OL�8{��oY7u=���^�'�G��xՇ���7��;�6��d(d=��������̃�8�|P�Q��^�f�)���HWs>߫��r>Ҹ�m����qBpCaG�Y�����"׸��r���n|�l��#��,6���^�z�]��5Y��K����es��)��	|U��D�����g��}9s���v��
�q�_Aү��Hb8��A�hE�2o:�� q��6�T/��n��*�9q��������7"�D^F��\N�.�/��%��k������7E�*�H�Op���fR�/@↥���"��fm.}��=�����C�Մ�k�A�M���V�v��sq�iV��}�V���[�+��"S��M�K���-�s9����p����'T~�&��C�s�ED����������W����%$Z^rʋ�wmk�A�q����}�*M!C������޹���Yd��++��Վ'p}����E�H�P)]�;E)w�	f��¶�*r V�_�Y�ev�8)��V�ㅯ�e��F���֕BG�JS��g��!y�q{���_	���xp�!nbmͺ�I��A�G����2*͘C,?M�7t[�Q�_Y��g���#�����\�z�"3�U�7��K�~ЖZ#`�Y�g�i�׳��^~ݦ%��:�=�6�EK��8ѻ�uDM#��F�&���K+�k���!�5m^W�j%�9q�������U5�f�L�0q��#��-������MS~ X��� S�t<)!=Ug8�!<�����4���HK�׺zO��0��Cl3PA[L2Y���VZC����C�c�xp:���-m��Ug�x
0�5�F�-H@ƃ7+��\!��6=�hm/�9��h�ϊb�u�K"G�8M�����2'L�T}�.��A;6�.n�a��,(O������X�H_�������p$�� mB�`Aw�Xg��m�Ut�go�x�>;ȗ{U�ז0�ô˰��-L��#y�˒7�C�)�`�`���F.)��y#m�{���� [c!q��\7 �)�Њ��`+]�N\����p"�����j�/���88��\])���2��Q���t�`�ko�`�i#O|�"��4����D�ۄMKrT��j�Q���K]?�%�RH���I����K�n�5l�h:��|C5�}	�l.���Ÿ��=���O��,8��AH�;������ma���5��<��	̋3X��(Ն �c��p�p�M�����ݗl��z��o��A���뾷�dX�����d�T�A����h��^�GOSx�4j���ށ8�CK��W^,��L���ǵ�7���!��w}��KP�L�Yӈ�7�ڑq[!FaqYd?�3[�v���t�Wɑ�$F}��:*֪;�?qB����]�ټG�fW�����Pe�jW���������k�N��,O�𶆠}%y�!�AR(��3�k7�%��ȑ��_�.��t$#�%H6�g7&��8(����ߧ��1�멯bwJ��X玨���cP�o�d�=Û=�CEӅV�Uv�䛹N?��K�C��<��b�y[�Y�5#�7 s4�g��{B�������P����z�V"�����Ҝƻg�ͫ1�=�����~t����XY�����t\�xGrR~�y�����c�ҷG#@/���^X�����`���[����+ʙ8���C��C+��E"\�8঳v�>'h���A��b�/��G,��E��Ň����X�I��.bǳM#�ܪYk�r1�u��u\���~d����K�m7��r�K=pQ(�Eu����rU%�D^d\�2�0[�:T������3�:C�&�d{���k@�j�S[ �'l�L�XQ�{w*滅�8ޠ��<�!�0��K�Mp�h`�4E<˒孨C����Zw������]��L'�k`�C�a��^t��ɀ%�1I���A�#VՌZ6�8�f����J����;��cj�Y�K��˿�/���Yw?��@$����SM8�6x_1e8����������/�(��Fֳ��m���}�">6�t�<�����II�]��,�*�*M�
�i�<EHu����{
�QNb��l�5|�{x�h����Q�0gK���®�c~G��8�VO�3Fo��}�6��ܯL�ނ��n��J��z�ʐ�Y��\�$H>����8�T�|I�Dfg̷?����eA�" ���\)O��C�,�c��e�ʸ!$���:Դa28/̍E����Y~J8��3"x��X���g֭�,I���-�ۓU>��t�7�b�K�|J�K=��J0Y Sk��n����D5����1ōk���7�A�u��S�����~��Tm�&��#��k�I(fՂ� keш�c �w K�w�Y)���p����2�9�:޹�!�v&6�*�=l)���8�v"&z(��ަ�Rҹ��,��Z��zx��ћ f�K�M[ַ�R����W�R��h����w��9�_O��H��!��c�1�ȄV'Y�i=O�µp�u��Ԩ�������;� O͠`��}0�Cf�VF m�������R�b�S�6^A����ǫIn#�?���dK�F���,kK��|5fY܌�������-�6�R�0/��]Z�	���RBu�� %�S�>��n鍉׏Żq���@<�L�r�0�y�g-���QUY���j�ԡ:z�s��A$7u�sx���q���-��ijl��,6�Mu�7��f6��֐͠ӏ��$ 1��R"�m�!�Գ��<oդ����\4����픍m�?uK�/�7-,'Aw�G���-���_��Xs� �<�C��U���D�2�Z�s膴}�e��l#yѷA�W%��&�ڪ��f�To�gT�Ȟ�F'���-"MH{lc�UΨu�C��)��H������� ^V�&�`MWQ8��Et�;����N����"[}|��ul���̴c���x�4zK��y�#�)����z|P� �v�v���9��}%<�2��r������D�����ǧ���j~����M�=f�\�+�'.&�[���ׅ�,�5�<N;�1wR�όA�����ϟ}���luKn��x�~�Z܋=b c���P�/��
xP齙Ș<����|7v���L��+k����)��ó��~	��Y�E�Ց\�8��@�%���i��X�ú\����K��jJ�*S Q̇�B��J�����*t�c��ə�|�aNA��>�ǱN�m)�����!��8�
��b��݊%���k�l���#���H��� �fT�	S��^-�Dp���e2v���n
 �(&t�Y�#4%FLtP��#<�dȚKQ�9\w���u���X���G�Z����|
��u����w1���m���@�ݪ��;��@[g;�Hj1�3�b��#i����1���,�`,,|�E4���wO�d��j�#��=}x�a�k��.�)5��<�W6����J�}ZJl������Hb 7j5zoդ�>�L�����FG[c	�yA<p{�t�H����J˓�_�͇��F%H1�ip���ɃS��ꂊ�"������t-���R�Ԅԫ�5Z��s�c
<��Fz�I�~���K����%�Lkk�}�����������Y-�f��ޣÝX8	"��~Y˴]�~��S��u����i~����t����KoFP��(n�+��շn�jD7Z8�oi����hn��BR~NA�t\9\�n�^��W\����E��Li���)�XԮ��^�ԍMH����Xa���b{n�s�3I���H�S	Iű@��f:��@���`�%7hv3֢�)o��qv�E���RF�9`%�Y�M1��7@;ܚԐ���Ur;����D%$���dH�J�F�d-~��>�!�u��P%k��#C���Nx�)���[Z�M��v��Y|,~=��SU��g���#�Th���6���f����U6e���m;@�`v��Y�̻^�X�n��y~�];&�˲��bAt�z�^*��Z'��`]��>u^�9x���\�r'P�����1�,� ·�wZg� ��&�Ê�|&�Ȓs���3���Y��2�x�w����u�	��j1�_C����tw����㦕!)�%¿6�F>��u�NIȐ$U���"�-/ף���
v#���K?=E�D��!+��q��c6y�p��;
 �Dy6@�7#�}���#���.#��:ݼ���Pe;y�4����$1v��/�����Y�`㩹(>>H1��	����q�;�	�?�ZdT�긯��]�������X�����$�j��Q	rg�@F�ݏ�z6��nRW��vLW��J���.��U'�E?��λR\Vn1��(Ũ3VB\�,�������W���Tk�������zu���Z�\\%�����R���.*��M�cV��!w���z)Y��ض���@�W2��󕕑���jj�o���1�R��&?|v�VN�>�LR=�Px)ZC��w�o��"Cu��}!.�|D�.��iv)E���P�C�8���H�a�l��Þ�A*:!����B�+�1�ky�]D� ���q���T�Nu��52���L���Y�E�!\ #==���/�C��) ��^4���V�����72�D�_??��
36��KÖ��לl��{`�)�yFfO�^�~������C"P��3�7���Z�hV$��R�;���fR�KK�3f2����;+̷#p�LEk��O�F��(�vs���0/�Z�����s���c��"+�;?����R����.as��jQ�M�[�nu�ؘ��>��Y��1檡?�����J��wd��O{�x��)�;;Ч��m��v�a�۴p'"�<�Zu����{aD��c�f28�����Ph��;'�̑׭�^CE�T���(ڿ���I%6�+yS��ܫ.u$�k~�sC!+����*����=��9��k�ꀚț]�G���yTX���o����J����6����	�JvFP�y�d�evz��D��a�O�S�D}my>[��ػ��\>�����o�8&e�����1JCW#$��m��@f�g�C�j�E��~��Ȋl��n4�Jqέ�ʨ�ɖɏ�sv��W��(N���~�۲ ��6vU��U P�*��O�ݎ�n��W�M��;fU�4�򥴛�kSM� ;,�H$��A�Ϧ��:z��c�e�5#���n;��i�0�=U�TM����u�s>WQ�R�jDI��*���`��i;�w[}�(pc�A��0jǅWuN�=�o��S+�I��͕��pn5�����,�w�e�82��>�AD%�$���n�9ѯ��w��� W0�X�-J�r���E�ًofe�7�Dv�[i��T��PX%��f�^]轛9D���Q�kb3��}�B5�߸�zV�m'<�҈�ߐ�ԟ���P$�\xt���2�J��!�,�#~CA}S�<\�����7{QC��&��5Nl�2�&z/��d�c���>�I�]�Iz]��(#7T ��e��[/*����#�oD���c��Jؗ,,/��|��8�+(37�%�%�Ԥ��Ÿѡ6a�v�eb�,*|pu�H�t�����᢬����K��j�(;ٸ�&-���NH�$�5S��+Q���������-��e@����J��VP�f��H$FBU���_�����{��3r���A�����KMw�֋�� ^ݧkU�-0vKeKH�l�Š�|x��sJ����ٶvbF&-�����4�e���N��1F���j���W��s_��a	T�p'@o�x@F�#uӞa���(h�jʺ�ax߹H��KRS0#A�7�Q�3��MS��_.��VD	H'���@]���\�ϴ ]U%z�ŵ�1�{f#U�A;9O�"��V�=b�g��K�c.��H{��?�!Qgg������x�ޮ�"�L�����MRh�K�_"he(DL���@����x0�..<���a�!� �`#CB�v@�o}�:?�xT���J�t�5�9<޲�U8��[�?u�R���|�Z��#��r�උK_z��(f��c��eSKo��֌�Β��h�y�,�����W/� !��(�2�������5�^<0�<8x:�L�_^m��f1-e��@�:���=���M�����nˑ�X�"lq1�Q�����4����ھ���Y��1G�LRM�f�#�ί���/��"��b����JV1!�7�YO!g� C�$�!҄w�u��(�2���1���D�:��/��I��d���d��������G�YR�����!�&R��:��G� �p�Z�}������tl)��#��]���{���H�E��?G��=E��|3?��2@��>*7��������v񬚯��Zu�O�������~FN�ne�!h�϶y� v�Gg%���l)Y�SK�U��mPO l��:'�����)���-��!RT�]O�o'�yw��f�/�Y��"��w��aP�{�*��r7�\��Hb��W���O����Ѻ���mx�+��R�A�e�@@%�6&��+#�0����a&���+?�]�����y=>b�]�f��\!�v>���V�E��Ky;c���9��[;A�7��j�i�X����(����\'��@�Q,�x��[�}���m�zx}	������|��7����X�l[~H��(�\5}�A������ڜ��h2;�rE��`��7�.���c�9���~�7�&�;���ᒀ�
�ɣ9.2�<�X8����o��%��_c�X��W A<���ԗ!{�ݍk�����C/��{��{� 8�{S_a{��}�u3�Y����x���!s��u�.P`_I�})����B�!?��'�n�ZK�m󉔌!�_A�>�cT2à}�O�b�݅�]ٳ�8�:k���G���S���+V��-!�w�j>�KYz��~�D_UEF�9�=�Ũ\Ԍ�'	��|a{]:�*B���.�J����-�74:�I  �W��س\O�D�5����b�r1��CUX�
v9p������re�&ޯ\���[�e�Y�*��[��P���q..?�����Lp� �Z�$�]rO����Ux˦k��'�!��rf}s�M$�§��K���v�Bq]-iGw�UG\0<x�����'��b�>I�"ށ��pُ������%()�����y�8a̯ 	�o��q�=Q�%��W��d�ϼ0�Pm�X���iw�=o������7}A�׭e�tf<��x�ly�-y遳t���Ǟ���8fh���`is�'�d0I��O���n�:���md�+��!|�u�eJm�Q�^�~(�YBoz�%y��Ǆ2�R�S �Ht%;��'[ŭ����u��'W����������-���b� ���,K��F���B�ꍠ�$F�U�����]�l�DԶc&x��S�C~�cB���	Dj�@yR~����G����62�Һ%Hƙ	U�-E,.u^�˓q�)��-�0+��3B�/'��t���vbDN^��DK
B��_���Kv�~h��RAb)� Ec��U����˂fRT��jZT�BI B0��QS�gN������!��9��@c��\ϓ�%��[}'��^pW�LKJW��l�����R6$�޹�bG���eՠ��d�_i��Ŵ��6e�$����6�0�l��������ݴ���b�B����9S��J�]��*�Y�i@!����IC�$$�J���\Q��0Ќn��g����Y,�~7�@'���W��hDY�"'�(N�OB�E=a�b"�~��N3ޠ������^T~��mh�)��0�h�i�M{�����ƨ��s�͚�߳�LtK륕4Lu>5���|-�f��wa,_VP���m�bBS�������Ks��������iJQu��J&��g���������!��V�z��!5@�>�M?�8=�#�w���*��ʳȪ��+�^G�`R3U���A��͗�Mߓ¾�2=��x��w�"�ZXG��l���v�+6�
w
���߫�h�<�����������^�B:]���G@%�ձy��#ظ�lN�例�b��j9�#E�EH@�̉�aݠ⾆?k��-����(���\�a�׎�d3&h��~8_�I�Z%=�З:H�u�%��w93�)�I��5���&H�x���?�!�~�Z���Lƣ,ĺ���������M�%x�]��"����W�1 5u�c��w�N��O[�;%*J{Js�Kqr��*g�I��8�0c��13��0|["*FG~��s
>�^�T�ElE����f�A��O~�A�Ǐd�i4��*5�e��*]�Y],z�6�?��+��{�	k�;�U�[L�$/B�_�۽�����IH��z*֠B��$�?N��ښ�F��<�@^C��G���8Q��L���͚n5�J�/�V�
������}�vǖ�2��!P��Ƒ������'��2;�!L�u�y��^ko��렄	��5�/Eb������q4���0���J�=�ѥ�< Au�WJ*a}!���v���QR?���:4��ob;�����X���)�􍼁r���!�����+v�CT�ú:�'�9�D��j��z�#��	8�7�J#=�IY�0D�/ߣ��e���liû>���ikr����J��}?�����ڒ#�~q�V����=��~�S�'���/��$�����Fe��-`;�Un��,��(��|���6=�U���-�>�#���P��&���d-�C�� ݿA`����s۲�󄁂A�u
�����FQN��5��Df��n�^�j�}�Kk,�Z�d`���p}��S�����Hl�`�x�~��N�a��u]9��5T�<��m����y��(�H6������_�����*��[zށO0h��W�ޡ ��-����Y4�s��+
���_��`��V���<3�����1�%���1��#���n�	��)7LzHJ��F�z>x�.غ&�e��O���]_�NM��r���u�&�"!sQ/Ⱥl�Vn�~/O��	c��~d,�aq��y�V~1p`��K���JH&�lqѵ$߳V	����48T"�ѥ:o��(�=���]����lj�_��V�G:=~sx�폹WatM��]��p(Av+�L~�����L/B53�5�������Y��b)ј�����K8�`����;PIPF��c��70�k��i���f$�hQQ��|�k��y�#��Z�be�@Ӈ� Y$�����l�P�����ڑ_�5� �1�S��"_�������R^AJ%;�Y���%WPP�@���%�)�'F-��a��6���q������'���2��*���,B+C7�iɱ�^��е�%W����P�,������%.���k�y,�G���w�k���������\V%���SM��M���癥n꯸��E0� n;B��RD��.xl�N���I��55 �-�����	N��Xk�����@ы��W�s"�_�|FF�8��x�Tf�"���:�>x9��p�44��tw����J���8�I��6�f2�t�6�*[>��E���yɞc�i|\�r�R���!M���2�jVzr6�D �ЂxX$�(;�Ó[v-��@�?�]��D���ʑ���KB	���1�˥;
=��<0� 9�`�������B����)�V�߁������[�6���L��#���	�kS����hƠ �н��]�;��g�oZZ��c^�y���s��|���Mȕ�C�'�]lYC�:�f��9��Z�a��جu_�
�i��@���N�>��K�޸��\��2-�*�����u��lpO�ݤ�P!�Y�C}�6.Y�-��^�Q�P���D���-�i,��P:8. �6��t��3[a@7"
�"��v�=�b<���LYwn~� S)Jm-���=�az)UJE�&��Fo�3�QR��[*7�æGK~*h@�ә��J��r��=2�b�:gȌ%�l�e[쯭3P":T����+e��j'w�y*<>�G�'<�Hb� �4B��}�`����ڦ�ދ���"Z.+��r�S�ڮ��W�g�-�����@�C�]	<��X���w~�닡Y��<������ݐs�Y���+���kC�Ƌ��Ձ��e��l��C���{�}�4J%G&���`���'�[����U���s�9�,T\�cl7@uųQ�թ8D"�m;\V_�I������^�@��+30�eB��jR�5�W]�3��?�t)���=��/oЍ��V~#�!?>�~����E�^��&� pg�������Qo��T�����;5[v��Z�y`2tfV�����m��4��m�$V�b���Lթ�#rWQ�������ѻ�b��êԁk��-%{���L��L׀�C�62�B���s�� ;.d���+�v%-��5��&�S��
r��{����;c�;���f���>�<�P�dn{�즟���U[����C2�'W窓(R�B4�棟�N#�1�0���6X��B����2��s�N�a�c�N~HT�z�/�%�A_p>�6�&��z�4>"�ϖsL}7���l�GJ�c��6.�R�K�
������UKUO�*6�gg�&߾���4�S$�][v�wj9Ns���y�Ѵ*�.��eWXg�(�r�u���w����٪�^�(��8�Ts�Z�hrL�]�K�3!u���wƧ�e���&=��S@�>�^�?�
�С3ҊW�M5C�A��Kdױ-ױ=����E:q�ՅP��Cș'̺%�����t����ǭɏ�^k�m@�;W�&����h8zIV����DI���/�w:1�k�A�=�;y}� �m�����m���ah��0�e����j����Z�-��*�+�G�(#��T�]��}G@�ܩn���@�b��r¦��:3\�=&�9�6�ᩋ(���X\u��Gc��r,��|���@pm�Ӌ���̈́�_d����U�m.�wO���#5.�E�;7�ރv!w�N�����?٘ ~���ĉ�g�:Ȉ,Z<{<<U�����~+�z�ph4b���`W,���Q��sc6�����R�+�yy�i̇�a��D���E}wM���r��mU���һ=��-�4
���Y���ƾˁʶ�Z�̗��&T��R+�+��Db���7��Q�p��͵卦'Ưt-�kf�	L|j���G�ڵ/�=�7<�af5�,=+d�a0	���OL����b��?�[K� ��	�|�ՈXK�/� I���ܡ�$�KD�D����[����+'�ѳ�zC]ȡ{�[\�t��v�
��4�s���r����}Xe��Z����;���?��3�cS����fc�Z6��$[9x�J=a���j����}��^�_>v�3��2���F/�a����߃�;':_��]�d�M�����sxmGVz~/xŋ��$x��Ht�x�@��$SM] ϱ	_#g]���-�݄x�]��3�c��9O~��C��t�RS�.���c �~g��i�GdQsdzM�_����ŗ�(����	��;\.z�3'�Z*��j.��cf!no?Cg �^=����*d��?Fg6϶��7��?ƌ�\f��p~�ҝ�=>z��|B0�8���k�E��
��W�����duV0 5�����Y�㦍<yt�I�ؠ�ƯƂ��Ѝ���<�L���׽�Q�/���� ����J�ĝ��5�]s�\���g���@��d��9���<!� x<�����9?o��D��O��S`��"����n=uE4*z���"����
�;Q��Գ�)�c�/������6�D�ok��ݡ�:ſ�o"Έ��_���I��=m���?pDG�.�@Y)�ȋ�Qw�<Ί~�]/�*�x��~��;���$Ezq���T�3t�}v�Z�Œ�p���rʌz�2}m����<��ao`�=[���A��M���}n�����$#��X
��(Fz����9$o�T&�qz���<�2������q��W� ���ى���uk�X�����/�LE������3GE���k	-�]`u����js���8}����c���rv~Ta�9AAsZ��3;3�ch�	�G@��o��(��=e���W"�%��z����N&�Fғ��?+�BW��^|�zQtoؠ
H�8��@L��t�:���>ʌ3 e���y}�\��Y�AH�uQ�_�a~.jqR?�J/����Z�gt��������������*�}������$��~*��_����(�f��rt�m�f;eN��ּ�|($Y�e����:���+���ڗ:����Z
z-������nr���������v��+�]��׃��Ҧ{� ���8� e��L�X��g(����&3 d��((d�wn�G������ފcΘ51�pV�Z�gM�~!�%%���X����# !H����(nX6�g_�=�rѣ��ɫ|g9�<l<!�0c��t�L����d'!��J��Dz�#�R-@R���H�ˉ���	�5���g,N�c������y�d��5=z��E����J&���p�ht���6.�����P�>V���p����A�:Z�+@�p�ߨ����Z��x�L]t��>a����^�R3e����K��nX<۾�%t?����$<[�\��l�ܸ���9���N�]1�s��/�vR�lJ��hR䇟y5(Z{��k��(���[�~.0����1&���(��Ђ2%nf<��(=��	�����Rs����s%Z�ʟ�y��v�bfS�i#I\��������%)��e!u�u��:�0q�&g�Uț󼲁��hÈ�6��b��љ��d���Z��[�L�B ��J�����nD��]Sik�TQ��u;*�^�T�9�'���4�1����X�*mz
���]��� �E�/�}�xeL]>z/�+��~'�2�g3<�9�	��X�����,���xݰ>ܩ-b�������iVy2#�|�L�	�r>ix^�y]Ď'+������e�b�w��yUb�-`��(<[G�V�~a���J-̛ݡ?�h4�2���aK'=��������z�<BZD&^9ԆҒ�,���^�5V2bLG��U��`+�lV��,���M��%?n+��l5��^z�5�`&C;_���|V�Zo	�^9+�
']��&~^{ c��CdY��;�m���9_;�6߸���v��ůE��UJa"��c�Ƌ]���y:߆R����G������]�2��׋�1'�S��ve5�ג�%���$���Z�l����wt:'��wӷ�U^LY�2�1�����%c�o~�����KTJ�@H��\�����+S{�S�q��n(8D˅��=�m����;8~ŋo�k���3��ٿ��Z������,�W4:	\���l�+�,d��xw5?�iN��L�uP�v�׽H8��dS��q�Ha�(_�1Y�`/V�c��ٷ�dཛྷ����-U���]X�Z^c�&�$�D���g���N��;�k2;�g�C�v����1t�O)i'�H䳹������.'�k߳d�oS}�P���h�������߸�	w�i��.��훢�:��������Og����:F/�b��3����;�nY_	�W�O��k�����P_ j�r��a��^(#R���۽*�l]���{�ʋ9XԆE{=�U�1��g�MX6a�v$C
���j� ��..�[�?m��Syz.�`��<�����v�ı��_�4��7YVk��a:.^����Q5�:�`$D��z����"VƊ�x�@����H��u7,Ғ|!Y��H4��4u<m��>+�qr�_���GÛ��9�M��R��_w;3!u6��qt��y��1����l�	�;�����oTs� }��g�ҥ�\m'NN��3�}{W%.�b��T��}y�ۆtW˅uA�F�+@ők�yƄh&��_}�i�-�&\�Ŗ�ᩚ7J�9��a+_�_�A�~H�+_���){~e�Ud�@���sh��G��c�Z��7�4���͝m[���-&M>����+���!��G	Q���8����P������W�٠�M�V�u�{Y<��x�f(��Ri�p���&HF�*BN��mY�dϠ2����LWJo#��/(}�7Y%e|��>�޵U�A�˱�C`W��8Jb�妕]MվR�{���b�j�Y ��Uu��.
oڻ~l�wf讶�$H�qR���_�t��U:K�,2I�^2��5%#zݛ_�w��;���� 1u����ק���!��a��g�[����x�g�o���S�l�	�1�>�YW'���yEt/zb��$���V��X
���ūe���q�f�)�󐓭�2g�S����;fW3����~;���ӥ�j�����8T��eW�>K89�h�,,�]^�~z^Vhc�Ӥ���j���~���0O�&[\�z�w0䦑w�E�t��"^�丆�oEd��Ju3!g+��.��qT���n���<��8�$���M���]�q=/���y�נ�� /�7VVΜ�3\S�¿�p@͝�	��X�Y*���H^q�9���۪�k�g�i����2�"�f�Yk+���]0V��tq�;~�����:��5��� a�;���	�J-W�N�Rz�v��1%-��ˬg�W��m�8��H1���{)(@[�)��'�C����k�"[��+�ϓ��p�;R���M����9/���J�/�J�b��a��YDN��}�p����>�}�$�/��Z0�������P5�p˞�z�?�x:�y�>5���%��h��q�+˛ �"ͧ�����W�7����Q�@�\©�r��/Wy��~8��+Wxwq2:�(�-G��G{~�`Ѧ������at{�,j�W_ξ\s�e���Դߚq�k@�+��m��VYm�������V��>=7�.���FD�杋"�x�d�z��q�
�ix�~�?���J��nm�:���>>
�xD%��~�CsZ�,������ߺׇ�_��k��}�hS.��=��?�/(b�j��j�����oQ}_�0~DAR�CBRB�[��Qi�N�.	���fTD�K�[ax����#���\�̜��ޫ��{�6�v.=z�s[	Pnx��fّ��eԓ+O�z��|y�����Vn��,b�<68�	���Ӗ�y�,��N��$9�/2���^h�)lyMA��!�YZ^��4{���o��x!e_kj2�B$��\��@�,q��W�}F�T4�4
0����@:���
���̽�;H�6y	��C1�����[�,���V��v���e�N8�	�$�~r�k�a�t.ޣ�.D�o�'ٯ�k�E[}]�lLIKWx!���7��,�m�g��6�q���eKNJ@�ڶT����-e)��_�a9�ec��>�_�g9����ǭ��#��u"�b3j���Z�wy��]ӊ�!�R�P�����;H���&�Cټ��D���V�Ǐ�ҙ�߄,�Cr����֜�� � 	���(���v��ʈ�����x�@γP�{}�K���%��up�U���1u�~E��~]yEq>&b���7�X��	T�1��s����z�W �6D�ܻ�&�ڞNPT��� �&/}n����h��dI8�lj���R�����Qo�7�cJ?�}I(�Z���<RG�6���,��}|Q}~��6td�p�+ްa���O�Z,��?��vpKE��m1A4ً�?D��u���o&�x�u�oW�Z��d�y���NC't����O��{y�놀�7�	��|��Q��{
Wz��(y��>l�h���4�C�	W��%��W�ټ:���6(�
�R���.D �ӼA���b�����F���a��/]p�)n$]�� ��s���H.oR���)��I�ab%$�XY��FHA}t���UD"��}��#����Ƿ����V��6���,���>M��4����\g5Z~	�����b��.)�^�u��C�e���9�|�c�ھ$	����K~�5�?\DRb�Ux_�_L�\��<k8#ҭz?�����g���q'$��UZ5�֊��f\{��YV�Ҡ���+��zA�kW{w'��8� ������I�.J�1_��x����Rb��6�ŝ���5P���<�c��c�I�lx��YA���8
A	��}孮����� -���K����<����������ڸM4�a�ĝ��GU���2.'�'-���6Z%�5뷘���u���m:?Ɋ9��T��M��}�U�k��)���'��� ����>v�Y?�V/\=[K����k��/sؖ�����áR
H�x1*���W6��uHV&�~�gF�(=%d�V�B��ֱy,QM�z�lܬ�@�3�W^>#��-Ց����,d��*���1�޾�ϲ¦nC<�kG<4���g_���Fٻ��7��`ߢj�=�r'��;��ӓ�54�}:�}*�'���!��j:�O�u~��{V��Z���^��lF#���&Xl6H�t���vJG
�2}��]2�E��k�qo���.�;��+2�1t�ZJM���9���x�r+�k� �߶NJ��G����k/ ���%S�_�p�=L`���
�k�TE!t\ZQ�5���X����Ԧ'�(JE��9`B��f��g��!V`�����x�5r�Y�����>�{�KK�NɄț��o_���&���+���䋾8���߳�
�0���Tj/�������8ƕTj��X`Ã
�ښ�~��m9��|sx]Z^�bdi�F�;
����鎭~G�O8����ӽ���]� ߫��=d*%�̇�篏;��������·	��7s����'����/�X˻O�M;v^�1�Z�}�>�w���BGNU�o���F�1�'���}�.���P�����0�ȰZ�q9���]|�mq2�"�ۊ�=vi�'��z<2�N�R��	Xtη�JC=����.��g�Xl9�u�����~8��g��S����.�o*E�C\��|�!?,jP�/f@c�(	�d#a]d�g��|d���y�&B� �ȷ�B֎����uNo�k����B��[7~*CJ�D��B�H{�'��B�|s���A�9�}�����������ү��+���8XX	��Jh���N�"�'v���+`X(��6�Z�����7&oL���ar?J�8Y{#��T�����q����c.j4#��<-�Tr]v�U�W�v�y��{�Mc�u�k �j䁢2�; �cT�OFK^(Y�g�c�ߛ[���`UNYߥK�P�zH�~~Oh�؋�l*�Z9�-�W�f٦��l[G����n]E{�ש�ZQ�K_�,j�_�^��&��]s�2@����p�] ��~��\vU��Q�FE�2c��hq*
��4(�B/w�໹�9H�|0�P�_6���/��?vsb~�"ٸ��y�AR�0a]9PT�.'3+K1�,����l�JxYy�+�O/ȏ�M���R������%we\��'��9��KS�{��gj���Q�>P?2�^��.V����̧��c��j��q$G���ݳ����Կ���^K����9,����BD�y�qAv���7(�K��� �F{eN�q���R�ph}�]�Q'�t���Bh8`��/;
��cX0��y�>"�.��/N՞e�n�/�q@P�V{��e���7��pA�Z�|ҏL�Z���
ꖽ���3�����+O���S>�Z{�3�%�@�(�r��Z�%��M9�kR�Ț����X���+�{�� �22�^��)���q�FΧ�z,�7sj�ص���`�flġ�ٻ��3{X�:��`��.)����ݴ��H����sq͏���M��6�����U��)��m���臆��ۨ���k�a��8�)�(u�K���k�+��]q�m����M��'��%���� ��N  [��+n�'���W�q�ĸ�4�n@ᮃ&�����Eb��o�A^��ק��!�:W��$��׫� �7�1sq�Uk��*�0��9Y��5���x�5z"a��+?�zls'��q�$����w�����.����JSd��V��'����^Mml�l6�᝔�\�����K�h����	ӆa �ЬjwӒ�4�J򕁼����I��a�µd����Eq�4�-�-�P�e��z0�WM�i1I#�v��5�R�37�Y��c�Z���,E8��h�t_Ք���������T�����?�6�j�j��sa7�! �aP*�˲�fd����IɷU�/���'��8���^�e�S���]-���$�S�m��ˮ�g����c����EdD%Ϋua���e�]EC�l�0�g�	��)��t0���q�bA<ϨRq��A�~�����s��"+F�[��8�A�����ϝo�o�C���؀������oj���GJ ^Թ9��Y�K^E��$���im��W����g�ie�3KD��m�7;J�K�/�V�y�����}@9ρ�b;+�������[k�B��0�m�ͱ�>�^��|�
v��m��m����v�*��vY��yq߳����l*W竊�F8 ��L��=fdZ���D���Rs��D�GX�:�2�7m�lx�B�UZ���y�m�*
[��"p�`Eq��*�\�p�����o&֤�o��Y6~k�W����5Ql�B�� r��*�u�������|o�˝�}���3��V�C�{�Q:��DZ�;DAɼ�+=	Lw��/{7a�$���s�j�]p�$�C+���z$��l��!C�]�Ўcv 0�7<X��e�s��Rx��I��f£��G%~���{/C,u��2���cfw�v�ÛSW�Sր�H��I���{��!��������s9a���[$p����gcs�=6Q��4A��}��JY���~�C�K�^<�/�j�[��o�W�?}�S{/�%���ݭ:�����,����,������|RU��@�)/�B����x������@�(e�Z��2�ɝ�%Rټ�����y�������'W��?�l��ڭ�i.�˼��������g�Ӯ=����aP1���Y:����711�����jU�L�Q��3ts�-=�>�M�N[�H��� W3��`���t L��4��7�ha��w��R誝��Gj�Ugٽ߸� /RZ�������$��B$�w�Ϋ`^-eW��0[�#)�rI5���:�'��PĒ�/,h�2��?��m(С��"�H������2Q�/�?/(+�$�ϤqgmT��ZO��[d 4�����ko��?CI�5k9��k�����>U#�m`��0���)x���֜m�����˲�wcu��o����B���a�f�x*v�:r��l�x8ܶ��k9"$�]��d��>�z[�����d��ɏ:sk�%.�MDn)?L��_]��C�)�%x���e#��$?�Z��=�覸o(Uk��#Vrx���'q��I�sf+0�>�,�PQ���NK�U�s=�Yz�G�I!���m�� �2b�Bu��!^{-h�����RG_E;�ƛ�~��'V��rL��+��"ǅ�B�Z��7�����ve���{-���U�TL�踄<C����=q�5�d�o�wCʀ���	X�
��?M�{;�e��G&U�惌�lt»,K�(���ۜ���O�.ǿ��=�%�e���)Z��6�ȗ�AE��ל��Mҧ�4�eө�ʊK�Z���"G�&7V��Ulp-�VK?>��6�a 1�&=��W�tGi_JN�J�8�*���h����{�[����Z�{��h�gKs.���9�����M�7���t��Ǻ�"A�s��<�>�# �����f���>2�e��}ѐ��]�3s�zf�!45���hk��}�ev��=���%9-2�����7����t=����
�]�s��7�y��A�C��� nR��+y�����T��'���?��^�گ�\����G\��}e��r��:/������'���?^�UG'�W���8��!L�Dȭm�r��7"h��yϽ��"����1G�S�m��ַAJZɽ�5�*�ҏ��x��2?����;��6��?������d��#����̥��N��#o��ULÒ�I���e��=�l �}�7��cxE��Y'U�D-7��ȑ�ܹ���#i��huE���3�o.C�m5$:W&6� ��`�FǄ�7g�;o&�~߻�g����#�nu1g1��9��׳�óf\-Q���ZS�-�O�(��I��r�$ɶ&״#�����G�-�O��h�i~�d�q��u������U�&eC�:(�PU�����
�7��h�=����jfi�A�R6��w����"�Ŏ@����� ������w���hj��~	�`]{V�����fY���P;Ho�(�MD���^�y����x���E��L�ܐ��S[�g⣀U��c�%��I�QOP��.��� �t$X���J�~a�Ns�_��ecv�%9��4?����9�B=�L�Y���NwG ܬ�Ś���6�U���?)SYA�W�W�t��Z��4���,TrHV�67��2Ә���+�w*�b�|I���dt��O핲(��@π���IoH�j�s�"��=vsp���i����D��-�����(�e s���	70�LLҹ�a���q�yc���G�j�j�l���&�X��xڟ�O�mU�w�-���^ �y��"_�(?�ęUH���TT)��SB�NDa�����!�ę����CBX�!�?�K5�Y��)�"�|iQ�E8&e���a�<���꜅3u��'�Æa��Vw�=��4�gY��yY� \����Ŋ6�7��☛�튡�U�r�V����ꍼ���U�[ƀyC��Q2�Ռ��װFK�#�}+- ���ꨠ�V�&(Em�^�\�y�����pSy� .��P���o�y"��ߕD��J��)vP�#� q?��=�Swh���%�xɬ������"���u����O�?�Og�V���ٔWEI�p���c�6���ۥ��Z_`�X��+�����Q�����T�s�ԟ�u�e�#i�����"z
���� *Y+8���!:���EBG��)����y\.��{�-��r�*M/!X���'ͮ=�r��Wl�Y�=D�_؎idv ��9����+�T�g��d_^�<��K�뿰?)f��\�|�ڣ���4{0%Q�$�'P�θ��ۏscVs�~~��n!HZ���q$@��1:T������2ETM��}���l�P�2H�Y~�[d�I$����>�H��1��'Z�G���>��L@�D��\�H�'��U�`g��IVWv�\ �`f�eѴg�\�qy����N������ழ%��W�U�%����5+X/���"v�_�iM��\�8�%�v7{������V����n�����I���y�E��h�^'�epy���@K^/�x|��w�}_�j��4�O��<�����4��T���&�˽)Y���$�����5͹��ʸ>qG(��L�.��5]�z�+z��Y=�Ƚh�ݪ�O���������E(kM�������p�X����Y�1�{bU:��d��D�m<=w�b�$��^=�S1OeN0E��^�����ܝu�K�m)H(���e&Kq� <_p����s�}Rp����߀{�Ҭ�P�{ں�eMn���rH�B�[c[	Yaq�Y��ˮ�n�}Pk����p�����>t`�v'?��[b����b��5�X�ښ+�n?-T�8싏��N�/��ϝ�|E���y~`����/�����i9��L�u���!,�ݶ����{��� �ԅŷ�V/����X+����oc��"��*Zp�$�i�f����Rr��^�Ҙ�U��I�ԯnː��8w9>c5=�댿f���aa�F���E2\��mʞz�yҶ�'`�*'�,�-���ES����=�~:r/,��0��m��zA 5��K	�p��5լ��H����Is.�nV���U�o5����)���l)�[�:����CR:�$u��y�j�ww���ٍ߆YiL/h,X��P���إs%=�H/�%"�0��W�v+_��|j���q��?�NQb�q���a��O��q^S��Gs-_Z,��*v5��mWD��N���FrAoM���|5�<�s�U�-�\����V��3]�V_�Ψ��}M܅�Cp�k���pcT,6ϨB�|�� �gO����ڦ�����J���C�$�������Q=wn�`1�ӆ誁z˰�}]����
	O������h0Q����	}/�M��*0[�����ǭ���(;��~ů��P	#�h�2)U��~���%�$�:̕�[e�G�S��U�z[.�IH��,�`�vdl1�.�yw�#E[�Bt� ��;�~�������6Yݸ�ŷN>���6�Ycð�s9_Ώߟt�^/Ո`��'�2_c�~�~�����=����)��<L�_����G����
Aq)љ4���^�!�!|N��qSx�"hl�)0˙~+Qb�f�!��١��NʑXW�6G�@LW��%��V�l ��}!C���Wi.��
��MtĊAl�a�ڱE��?/	�x� �LP���?�@�{߅�[��z��z<�8��N����ߒ,��)����T-����.�������}��h�luo�C1����K�ɼ䠩@'����D�m8S��z��Q�M���'�_�����K�Ћ4�J�Xq�h�qc���Տa>g�]U�'����V��C@���K�We�jأ��g��/���[iN���8�+1����*����[���Lb/��%"��o�V~�%|��Kv�Z�+�j����Վ:p�;26��#�*�t�U�h�)a��:E:��^\����O��[�;F��뢽��R}*d���/�XY\��琦z�&��D܋#ɘ���FL��J�>�N*�r3;,�����p�&����v��{���
m�m���Z�O&|Co>¯�M��$JY}��b���4�^ڑ��;XNc�����#�Qf͟}����:��]�0���ӣ�'��K���%JT�@d� ÔwO���� %�+&�T;��Ì�
�7�͸�F�ئs��/��o������C�L�a��rÛf!z .�V	��p���ʒ�T۝q0���d� ^9
P!g]B:�H!��9�w٩D0���ɔ�F�S���~gx[�w��$���RIP�/� x羁m���� �B�W�(�k�(]!U="Y�� �s�|g�*hwynܯ�|�vqy"r�M�K�E��A��Xvʔ�o���'R��b�@��+|1�s���X���wNQ�jM�G�$j��σ�Zv����^ϻ�2Ӏ��r�0��_�_�~��آ�-��N�kY/;�^Ԯ�R:��'���6h����(2Z�"��	�2핊�qi�_�=���>U�������tŪMx�T=.��)!�5$~��Eز�J)�Ŀ�"�I�ؽ�!�>�D��팗���y�Q<#ܺ�a
s�y�;�G��{0�"Cd޻\<nz}A��gw��\V��@��k�7��Vw��T?�+l2&���&�����b�.��gL�!=���f�)l9�i��`�Wj\g�^����!��.vlY�E�rI�}����+�Z���;�

�j˨�G�{e=hƄCO�N���PmV#%�̈́~���z��L$�{D�h?Fo��C��o]t:�J���nT��/�S�?��/���IX&�g=Y�q��������WD�g%�!��SE�I�4n��]��{������$�-aX�j���Raj��-�,��7�=�M����/!�����߳���RCb��.훑Gp����ڼj�pZ"=<�����,$���X%`Sx>��,��J%��tI�Jk�jOA�*�+�a��~��������I�g2.V�������"��Y(|��G��YX�1�Y$��6%�� �ᘘP)���wD��,I���s)���t�	zy���X}�k�t2�����v�#����}
����c�\�7к�$�؋�������P�]�.�k��_���n�/���Ɔ4��n4��@�}c��Ξ|�B��Ȑ�\�6�W7�C�� Yݏ�YV�P*��.(5�=([����� �*�Z��R}��F��M�
�fR�o�YrU�T�d��*.��č�Y�ώU�Ba����7MM0M9{�&������߅�_0Ξ���z���ͬP~A�S�@n���Ѝi(��0�#��͚�38W����������^��x��M�}96<C�&���̿��u�R��s��v�bl�=��Ci8����<Y�����_������Ҳ֪�H������9�PI��_]��	U�P3������#�bd��;ل�0�U�vZ+�y�`\��"s�+�:��\� ?M�/;��g�}��uj�?�J�����	c�o[�6�����Rݓذc��g��#'��ZVCD�5�������z��w�\xT7��G��֮���g�
��D4i���^f�y�_��1�m��+S}��O��ď�u��ͣA}�>��"�&����_���$��M���6��q߳#��>����o��ڿ��b�%��S�Ѥ���L���ي�#د�R}r���H��x�k�턝'�2c���X��zY�o|��G�o��H}qʱ7�)���_
�<�hdl}��kr�݁m��U��9u�g�r}˜�aՏ�
k�Y��$�;��~�UtK�Vo�~�n��Brx�E���Vw=r�<�#�=^I�c��|�](C���d��!��k��"���FnKw��CDUh�J٭�q[���'c-�~%���}�5��1�P�WZ�Mg}��d~�O��z>���#{{;+�Dɠ��q��w�������C��R�Yd��v����>E�c�c������H�}�Ǉ�|KZ�yv���>}.E'K��.c�T�J�[��>u�)@E�<�����O�\�-���o?M��g"�}��p��et��R���nX�!�Đ��;�Sh>�+]�x�ق��)��%w�iS����k.��g�-Sf�T�`#��l��,�vH�o�o�"��%�2��eI�ؐW�N��P�0�F��gC�щ^���̋�*�,>�Q�Y�$�
x�[ϐS��x��6��|�:�'�L���j?�L��.�i�j=y͠$=}�

b|��Wo®kVu�q}��P���~h\�2�-��B��4Mt�65TR�&�9yg^�,��J��������s2�WR�k~�|�ƾ�bxl#�ϋ�w�>fe�r��e} $���3O��uR�P���W8o��r��^��~-U�)�t�Ѻ�7Co���� �F��Y�0�v��oQ\�À��J���\'`���F�l����_�BgY���%s*g^֪lWgW�ífW��$�ʖNasZ���N���a��Q��.��y%�[�Mf~C�9�LG4���z!k��o$�2ha�>�D�����H��]�������^,_&S��ƣu?z���ڭ�_������l>y���ɬ����y����_qm�c���ɝ	��Ӽ+���|��z3&�N(QʴIL_�?E#�BD�O�AX@T2~�*l�\���P��׮&��5��DKQ�#� ��ӓ�7|P5���dc��؋�a�P��'O\E�yą��9[f1�8��)E�9�s�Ǡ���>�4��M��m�l�rì�C�&���n=ٲ}^���S���D���Z�O�u�82��_����
?�������C�^��|�2O�U��Aj���ѣ������M~��Ƕc��w�j���	x������6�:�X�3�^B�4�I	�4�F��K{�a��9���_1�$�(�%�t�a�|g��-��/���4Q\C^�]����h̫<�����R)騬gG:�������v��-?C_�b��U]��t2�3km��Q�.�%��)�Se.}׊�Ͳ�%Z}��ǲ�䮡,wZ|g�14����Xe���Ϗ�}�ܵ��v��+�|��w�d���9�+	�x��p\���t��2:xl�ְ�����7��UZ��V
�����Z?Ʌg$�(�$�Մ
�ց�hb�鄪�ԇ�M6��Ұ����%�݂��Í+�4��������Oߡ�U�����g8x��X��M8M����'ѯ{��b/,�7����'��y}�2+�\��@h`$��m%�d���Z��_|�v�5D�9{������\@��e�ݦ~gq� B��D<t�c����%�^{r���zRCC*��|�N�{�ɜ�J�p,����y.�y���'u��B]V?C��uc[� 397���&,:�����{~���c$w����!��^:|��~i�J���R�UC��]Yʇ[WdMȇ%�MڮG)�O��v>���|(*EMzv��*��
����O��f�Z����P�xo�3�WE��mC�Ry>;ޚ}*���a�y�ʧ~�@U5r�|�	d�k�P���g���v+1�o��OP�MC�a��3)�5.�;���J+�g�`�����.�/�!O�q��f)%9,m�{Y��/����=%r��<��-p}Z��}�Ta��E�^K�m�A�����e�޲T��]��y�VZ��e1gf���� ���h�I���`�|ڐ/�ҽs���v��h�"_t���&��� �"��cE��`���u�����NM֦ͧQ��ĉ�/�y�į�����3��B�zA6��#��#W�ޅ<Ȣ�/53��;�e L����78V�}7J����E��iO��t]˞A��Uxr�.�M�e0�k�[��ŝ��o�O�H~�F��ߋ�E�?���f}U�\D���f]I騌�f�$�ټ�r/Q)?�9mB�)�J��#�7����x��]���vbX��{8����^���'Pܻ2�{�j�7y�E�@���.VUC��tm�6?�������t��j��䇍.���2B�c�Z^��Sxø���R2�����$[>�#��r��W6���q�3����Ӳ)e���i 9���_� Cִ���.�H+B�)�c�K�~" .]��|��#�c�fiv�!����+)����Jd1߃d	�,%\��r������#��������m$��Ip�qH牬���H�q�E�i�<������K�K�:�虸��g����a^�Ņ��%�b/�?:NU�h�ݧw������U�Y��j��N$��e�w�/���ֱ���Vt"��O;3.W)�R��>c1aq<�3�^=�vE�AN׬ѕ
�^`�/���2Bf�	v�9$���-R������WHQ��J^O�e�s,8��9g{�$�.W�|��zXNV	���
N�+�:!l1���@Q�VC6L브�t��Ġ-�&6;����z:�_	���͍�-ux|1v��~��:���%��\�1P�@@nx�L����Qi�ak�|e!�X'�O������!�&�\˻\��kr�(J�E�Z��E��=ԃ_�_^H�Z=m�7����[����0�@��15`V)����m$��Ij�I�l��0�S��+��gE��]
d� \|�0�8
��� �zc	
m��<�͉��a�<zх����X�=�{����z<�������}%���ş�3��^�E��Y��|$��w���tL�s�]�)�	�~ps�9r��)��f��׮��aE��K��̩�fra[��2��Ϩ�[߷��a�b$�=ŲV�����3{i�7}�=�����ڟb�C ��#����1f���E<�>�>S�\�JQc.�t�Ӧ�ŪO��V�S�bl��;�o;&��.�\:^:E�Hcc��)hnPָ�T�>�r��=-r(��e�� Q�cB���H�k�p�P�i�UcL9��K�w#zS�K�_� ��T�eg,,՛z'�ej4� Txe ������Dw"<�7��3�%'_� `n�����hy�Hg�xe���i����c�aΊ�8VO�e�m����ȁ�#��?6��Ke{�h}J��. Wy�������bL���8顖����t.ꕟ&�e��
� ᥚ�a��i�����)�
�(�j�cO�۳���N.S<�m�32n�l�)�0�o�JͶZmtx��Z���t�ֿ����,)���t\�����C��'%��(�&�2�������ң�67����]W�ޓ�mtJ)�st24I:�7p�7kLdk��t$������R�"�l��x~{,�����?���d���/>�M>v��x?��%���?��C߶\/�B7O���+�f������oX��w�R9�y����:�Oרq��l4˻f@�b����qE�~���zy����F���������<�G����J����J��������ր4��C�k2T��/̽+~��a�Z��ͥ��<��0�� r�P���R�zl���U��.w��&��U#(">q��+�[�Mś�b|=(��h�)�%Ҫ3���	!�L��[�UMQbq������	��7~�:�^���~��o/ B����<��7�%��f!��5��������� ���1�wv��O|}�$� �Wץ�b�7�!���Uy��{�'�R1�&����)����EC�8c�����ݻ��j��e���wDRT)�8�X7":sQ}Ku�m�bk)���h
~O�I!�C�Y���7���ϴ|������T�:��.s�Г��*o�������{�~��9c5�}�bS����~s��ϘT��]| j$ށ�u����K��Jw���gÛŦ[O�H�v�Y4ލ�M��ƞ�������XԴ�%�L��xs��7��h��~�������2]E�sб���H�����<�ZP��z��ڃ#�;XQ��Mm>�0�nʾ|"�UO$(��j�>�1�n�~<{3������[���o����E��/�(�j�����}��̤1���	#2���0D}�PuzW���dӶ���͔m�`�L��l�`]�`]kgBi�ħ΄O��/�܊�\�n)�(����I�~�ǈƨA����ќ>����ur�ێ�ے9j�^���a�����q��R@Ӛ���gؗIx-�:]ERr�D�"��o�����5~L��*�]\����;�j���rfMe�:/9�����$�y=8���A��L���@SW��}r�(�;�Vо)�LC_���bhZݨ<i*a-!@9A4yỆ���n��E��6E��Eܟ��\8P� �bB;��\��+J�u�������ϯ)��~o�./���n�����q�`��e!R�7q0J���J�>���b��)���1p�˙
k�.�$j�;ܚv6�#�#δ��8��A�V�~_V�j��9KЏ�fo.�����]-���Y=�����·�@���@t]X�)Nd�UO��+���k��"U��|'=�"o[�쌭��� z��8s�yZ,�,�2K�Z.��!bU�v��G�J��\��~3^��6�v���� ݦCe�8��d��|��,�ܱ1�}��V�16:uJ ɋ���R3\ڼ��� �T�k*��#�r/��un�f>�������q�z���K����떦*[X��.+�Td3g�QM��-�ι����F�A)���*b�s܀^[�Yr�[�� R���4JG��jȧ����V3�rBśf���iF">"xWN(3��FJL��� S�F>��p��Rv�X�--��}���z	�E�1�������M�!�J���A�d�r
Hf�&ᜱFn�<�Ov��+�eNCs��u.���F��7U��d	`��	�ciE���3�ܵ��θ�_2�(~ù7�V�ث�T��یÂf�����y�L�o�q�~s������2b�C��S߼�2��Qm���r�I��B"��*����j�6�>�`���3��+�#�������y�Ͼ]r�S,�mln�7�qҞ�QO+D">�s^���1���7=��&���Rۼ,exE�0���`+s��]��0�L�B�~k+)ٳ?C�,.(����y�G)J�	m�z�������ە�c_��a�ةF{�:;�ՠ�ɯ�Z�B��˅%����T��
O�' R�{^�O�	�}�|��c�kn�jP��=���=]��3Zo�є�ٛ����-ʭղ,���Q�n����h,\^-;�b���{R/N��e�t� 6(I���jr{x��4S7�hRS��R���ЍĒ��P��n�f��`�d�I�W^,E�Yoz�'Ku�W��Jy0V��̇���Z0W�ɸ�6�Z��h�&`�2?���\��fɾ�iO؆H�J��K�ZrT��Έ����g�$3��ʅq���A�������?���j0wSxQ]�e��j.a���$�8�QSVZ1�쌟�6O�o�����η�)�)Ta%�&!&Q�~�w(���]E�[���FVR�����i��g�!�O;�.Ց�+�C1q�L��yV>�@���&�Q�>^��A���DS��-+��Ɨ��փ׊}֞m_�4�����l[��8ܧ6$,�A��R�K����$��,n��/f_x3m�-�2�هx�c$|&*��_q�	7'7�Υժ�Q*Ӏş��@����(�?7_�O�����>��K��}H(u��&H+y��T|���z���� �sOſ��o����5�Ui^48o��r޲���l1�<+vt�/���V�؉������/G6m.���\$�튌�b��H�;�2�_�.��@u�X�_������,]���.m�Ӫ���Q��,���Y���tH����u�'[��-�'U잏QC#W{wD�kO��6�L�j���4��e~oK�|��0q��=� ��(����Ϭ��$Is�M����_�h�/���#`zG�� wgs��������Bt�]>�"�������Tf3�h:�
�� 1�fx�o~��%4�7g@���Ԑ4y�L :Ϲ�T�WW��q���Q�c�T��ь��D�)��G��b�����|Rc)1J�ч�^��Xm�	�&�6'��@;��*��i�����P%miŐ��7p�A�4�)������=p�b�e(A��	իJ� ��� F���Oq7wk3���} �Xm�T��j�=�s�#&b㧼��7����.W�c$H"�r1��;#�s�c���̷G[������ס�۱V�j�U�/3b�jԣB�.�o~��K !� B~���ʤ_Z]�k;*���-f��#�wV���ۇ��A�vw�~t;:T�LX/�U�a� ���������qj��Y�Re��H\k�+%��^.�6\�θdj�e{,���)�a��n(N�7�#A�W|&�S����̞�˫!���&c ��|jwqCP��%�E2Ѯ.Zn{&fV<6���,���I1�f�S��|�dcёfR����^�U��.C3�v�Q	�r(����++�:v��Z��NҀ��È_�H�ʚ��`h�(}�U��O�	���i6O��T�B�$��l�+�8�L�?�=.Nv�i�����@�,����{�J���W0�I�C~7I-�J�m����{�H�f�1�Q+���o�[h�}��a�;~X��'��I�X��7��x�OR/���P���p�#�+�&xz�_FϢ�gC�/$U���V&;�q>Y�m��G~1��z=�PHb􊪖ߣx�f�\\�6���}����h�k:W��WRu&{ E��,�L�P�BJG��Z-w)و�����	yH^~7o9T`���0�FRǑ�&������^�Ayw��Ҹ��n�3�����uhJb�7��lNKw���[�z	�J}�r��e�����w'��;/`[YXMnt]�\���;��X��=1f����{ؿ˚�6�5u9�	��)_!���L3�uF�ܟb�E�B���9��.�Ec����E*��=��.�cx�7hk�9�z%��a�]��<�ŭ�w���=�Nw�؎���6q+بx�՛z'JR=�D� 7T�X�.4����E�KcҒv�<����| ��	o��צ�:�2j�f�4�]k�N~���F��$��Xr�i�`�a�c˲��D=N]�ߎߗoT��i�ȴ9�4]uT�[�G���Wa@�[j(�n�i�zD����n�.)i�n�b�����~����>{��s�8�L�?��ն��Ou��ԣ�Ӳ!�
����ĕ�3��9ᵹx4S
w��d˸ִ��6�Typ
ù{��֛xu�U����D%/2�<=K��a/�P���XsM�,���,��.��#,�G�.kkm�����\�.=o����Ħ�+�/�?�k/��
��<s�p�ͩ��Q�:)� ��
�g�E~�"���q>1y\4X�l�4�]���&6�}b���kY�9�i��| �T��@^%��d�:�ɢO���őSk�%}T��vm�� ]�`�ĒcC��qW{�# �޶�Hh\
X%5ݛ.�f�L��?�qJ���A�j��.g��& ^��^�m*:�܎��iz0yv��!�)���� ������{0�,
���l��{ ���*���$���4�j������2�=��ǴL�I�%�Mn��m-5/�߮[62љ��O��O�.����[0ػY3l��N(@$�5)�R���fJ�N�����v �㺜�o�r�X�UU�/Jv�p�\W!�o����I�M�RiF�'	r*	%�ƹ�Mq�u��Sl���sz���<FK���Z2w�STR�]��J�Te-��
��u�6�՚��Si�Mn�mn�5�2�9�	���@�u�Y��u�2����Q_���XL�N��?Z�w�1#ں��|�"jUb@��^u��݉��֓*�>1����Hc}n���V,1(�)�b��A��\�Y�Q�4���+�c�VD����߸!)��Т�|o>e�}�Ձ�0'>�<�V��+j�QS���8.����:�5{-�qġx$�]\#�H�NBt��W�O�f^xpW��e����`u��:�_OjDEG�G�0_ԇ�#�1
�h-+���2�Z=&bXl��kp� 2~5�8�|��A�L��;`�	i���:{W7��0,:�QMcy�!�w�Ux� Q v��g�WdP��]�\�o)[��f;��_�F~�0��L)�k4�>�����v�?"y�����s`�g�FVՅ�-W�!lSs%3��6t�#;��òF֫1X?�׊M�f]9\V�Y�c��M>����>��Ͻ&�sG����j:��2�LZȾh�Q\U2̢$I@�[|Y4S<7���^��<����0�"1۴��P�e�{��E���*�*�X�����ֵdG�	~T?�ʦ�es[���,���QC�G9|��T��OF���z��*(���@�z��y�1�K��JV�f����}M���aq�u�����s����K~�S��u��tQ��N�#p�`�ꊍ������֬�ƬH�Q���ܫV�5q];����2�}r�)5-Gp�Ǟ2�Fث����WiW[��v\[{n����!cW��ne-kQ&�^�l�&ҭu�s��ð�E����U\�n{��,3�t��"�L.�Ȧcd����u׊�<{���<!��i�l{�E�;δԷ�B��?����EPR��i%���X;���~S��m�.�����B�6��E���L�V P��H,�x �#��A]t��Ia�amK����Q=�R�`��U6�S��N����N2�0ٺn��~�������\�]|��ď�Kl�Մp�A"5$��.Iof��'�R\�F��+w�6��ɓGbڵl�����P����it�n"��Y���dvq�p�9^+1g�4������{��X���:�Z����M
�ޑ�P�?�ݸ�j��Iv'$�ݮB����&�%�k��|��GLVt8M�=&V���Dz��68#
Xu`1~��}��b��`!���=�k�'QF�gF�[LU�/��NH�f2��c�?n���n��|]��Zp�_Xc�I{� {�Xf�K�9�x�_)��;4y�M.lk�e��RT�J,�����Xq��`͛;�O�&�U��*��d�}�?:�PY��/Fw�q��,0sK�a��6Y��N�WT;׌��i�:������磑i�GSgA�w��u�zfX���Z	yF	T���qn�f��n��[ �`��{��#f��e~g�mns�)=Q¿ ����UJ��iy����b �#�S�{�5B��ב/�K�b<�#��N3'PpY��|��^�����էX�?������R�1!\�e�?8��[�ãUD�7�C#�9��N�<r>��g�8����	��m�M�;�^��;4�KW�����t^G�����B�9��-[ܑ���BX�7
���u@H��\��u76�3\^���zh���o9+ٹ�ڸjՅ�w	7�{@8̾��~�g�U|r�kW�t+��6��i�k||ԥ��yQl�*3'�i+H�8x��w+m%�����:����!�7�K�v}�o���3N ���[=��L��Xr��*q���D�B�w9Lkx1&��rZ�����-�Y�G}+�)��!��X�5��Ĕn
��-����M������|=؊B�Q@�ݣ�t'�g��c�n��*��G�@�L2q�2x���UZ�H����>I�#>nmS��@����X�y�K���Ψ����I�wף,ԍ`�@50�M�3�i���I�l��-�K�@�4O�_[�>���	ި� M3����~��`�e���X�f�P�i���y��R�7ЌJ*�nb JM��D��:	<�~=@�R|�je�X0����� ze����-Z@�2��H1��2}�H*�������O�f��b���Vi;�h�-ǧ����G��h�dD�����5�����e�)hYG���)�p���cU�@����=�M��RQ���h�O�z����դ��ë��R;��_sl��:fZ"�DB�7������@�`SK����M�_���
;���'��]TG����2LQ����3�G���Op�65a	��'O��ܹ��O���L����M^�<9��q�τ���V߽V��kɕ�����aF�V�������*4IR$�İ!�;�m� }��f�;�Ԡ�R�LEbB����1._K>LB�>�b�]�>��T���N|x��w9��b�MR�Y�t�_'��ׯ��߻�{�{���_5���k�VWM����4r�J��jqS3�ȫ��mhK��&涤9J�qh��e���e�	�FFםS�����)�C9�\���=G���R����O��S��5��[�i����U��'Xx�z"�#���'�.kl������q>���Ա�tN��^��0�^�Xu9�9	<r�2}�Q/��^.F�0�^���aBq�̒>��~�+Y�/C50�X���^w�Y���ZF٥���<�ux��es�����^�~��Rn�ԍ�����%��O`!���	�C�`u���mĊ�;����� z|�����h؞�Q��m7������d�>if�.D?q��P��_Vg%�ї����L���w�W����T}9 ���rem؟>�s9)[[4���T��!F5��f$�D�!�Lq�E����kb��(�lM�@q[�Y�:y�X��!��Q�HӠq�7P����1�������߾�����:;g~=���=	&�������1�޶m���:=B�a�*���0q���.��/c|d!,�?�$���u�t��;˖�bE�vh
���OP�Nk����~^������D�Ҟ뀼�:QM�yn�l�����������n�t�C���G7�T��0�7�&d�4/;'��Q{duqj(�{�2=�`+��E-��
{äM_��g��t��u��MYsMn^���q�8��C�w��9��#��xU�j�nJ+�G�S�	>��D(��֗`˼��]��5:T���>S=�#����z+�k�-8�=]�Ⱦ(�[�I@���7�Wa�$�u��R��+�y�r��^�A�'�dPeٖ>r����Y]ZF�)�{ݬc4�v��5ݱծ�D���1Z��v�L���8����2�^���Y��#�(>w�L��u��_К�<3�0�d����c��������-��J mv���	��u�j��r��vb�-�;[�:A��&���n`��'hD��o�:m�w԰Â�v�tȫ�lKt�{���+�S	4��p<����9�{5��?0��<��Ct�K���M'uΣ�rI����r5(J��!���3�����F@��,�?�'L���Q�#A]��I�,��6X���^)�W�����%���ߌU�����	*�E!ĉ���K�6o�!�3r�	oM�ܯ�aE�_�C� CA�X������	�Z�:���}������v�7�xWy}��$A]��=�>�<���7I�4��b}`ޭ����ȱ�oßfn��u���ү&�TE��[�ɿT��[ǅ�\.��ه��whᨭ:]��Ձ���^���h�b��0��o�����]�3;@��˜�uU��c�������l�]�'5m��DЦRǋ`�~�r�k��ճ���v �|��f�Z����z�W��>=�����>��
N�gS ��n��M/��#;��"NE��y����/����\\c��sZ�?<��f�?����KȠ>�C��R"kr2��^ܓ���f��[=��7�A"}�<�N�iޡ1����.�[����Ab�_Ի��7!��`�fj��Ѳd'���Wp0?��Q������Y��ٵ!cwi�#kMM����-�K�{�d�����Y�1%V5L�ȉMsޤ��� ��i�-(�W�Ӎ�=�GND(}mvV�I���^�߅�\�N�t�%��T�G*J�G��oe,�s"�+0r��y>�d�U��� 5��J��Ò%է�.~��6��ƙ�WߕMr��W�o�9��R����O��g��e����s�������>�I�Fq�?6��U�|.۝3͘oB��l��dk^����sR!k��vK��4A��
_{���'-+��J��r�k�qS�`��9��f�u{#\�VV���@v��0��{׸���4�O;ФQN�  �&���@�V݀5U-��r�4����\S��?�6\U@HaCwb֖�Q�sr�X��:�|0V�N�*l%حi#��-���z�߮g@к�S�D���/N泶�ٲdU�z�:Au(���(R�9�6����k�tcZ3�����m��Uy����'��U�+�?�	�	��I��3�Z5��
�t`p�r�$
e��;���7^W���Y�z�v�8������D�-!���۶��,�3���m̚��A����Hw���[����7�6�u��}:ͫ1��U�"U�Ȑ�"O��Ӟgx>����H(��jx���y����ٽ4\tªh/�D���M��������OWfV\fz�.��.�Sir�Q�o�x�c:&4��僿^��JUuC�|WC�����f�bx�c!s{�X��m���Ġx��m侘Ԉ���9r����p���<ƿ���b���(�
��Yi����S�����M����s�(�h;��s�i&6!�g��J�	mŚ�_�S�Jq���  �[Ti���`	�zHb�����/]gl�����}����o\��6���O����-�=$}�~�&X��&h;�J�x�a6L���+�l�-�7f�C�}8X������E����9V�E[�o�͵-ZI!G
� C�ri��)�%=��g�NY�c_����(�_&���ąuK\[Zё�G7z(���l1/�MD��6���O	��QL���<��/��Q����P���?�r^���%"�,���k�n��e����T�,Ǯ��Y#�-�/��O>��X�������f"��Ѽ�ˡe�c�N�b�5���詖!�	�����ΰ�j�2}��n�Y��^da����}>Zՙ��n�B��-?.�M�~p�j8���0���'��\��>� Lc	H�ߥM�k=pC���eb�?72`�ݡs՞��3��:���|'d���610���e��e��$1�dO7��]p�4,�X`�?u�SB�1�̗y��I2<u�� �$L{c�r,����ݧ�����?����g	���}�(U�O|��o܍0bzǗ�X��1 ��5c���+�C��"��y`��Ud�y�Q���uK9��i��E
4cV��-����u�%�����n�E����δ�ؖ�̀����5 �ц��K
k�,Hm�v�,90.�� )���k^��1�{'z
o���m�Ĉ�U��ڝ�E,�
f� ��Ai\���v�J/M�y�fR����<n�;�>-��	W�`. ޯV�r����c��-�b'��]����c���N�%��E���U�ٷ3t6[�\�����@^�������f˘o3�M�bz��m����S�yrX����/1(-Sl+��c�/K�!H��X�����T1%�I(�NB���-/�ǐ�^6I��^�����v.Jli���Fn�xpS�zQ+Y�Q����M
�-Ŕ�+=��eIF�(�<��@��@�+{�F�;�����&!�vKh�B*5�������*#8|8e���i�:�*��z5�����v�������,�|�Z���6<���j�>'�m]+cڊЊ�� Ȁ��c5@����)�^�������f�ʟFO���U�� ��J�
i�
�\��
>B��k��-~a2Y�V���4�V�lQ_j������h.1��g����K� �qbF����l�h�����F��~��̋�vOi�x�y��2=�X�S�e�;u\�,�vb8!|�۳ X����e=u�y��l�d����f���Qn��#�u��iI��o����zo�5������.䪒+��
(ݤ�����W�8�3X7 ���?W�LJy��bh�K�K�yl#_�/? ��s�x��m�f�ήIʝ�zuW:Ќ@/L�����w���7���{���|i��B��� IS!Tkp��@j��G*��B�Q���!�h�@Y�n�sp	����~�����<����7U�Q�X��&�<t��p�|_�|�$���������7Y?���\���tq*�Ck�'�6,w[Oxz~6���-�S���m��?��M⽲�z���N��v��,9�8�Y�#�pc� ���j�MaB��˺�Ea~��RѤ�6�1ۺ��+�!�R,}9�W��Q6�b����:3S�gׅ�Q�Ħun>d�᳿b�-���m��(���a��&[�h��{u�|�iu�r&NI�m2����M%%*�^�Y��U��$�RXZ��L��믦�Lۚ�X�Hs w!	����$�y��n#I��������?�yn�U�UY淎ZM�n�0GݯE����(*�1q)|��E9��_%)=�Nh���c�0��t7��������0[Ѹ��+��:0���/�`����ca��Cg���9����q9��5��Z�i>���6r��2H:@! a�~��#)Ҿ�}��-��7
��չ7��x�ֆB�½������TN �{TK+�����t�Y�S�2��c����7��9cƭU�B\��v��LW�h|�]ow���y
�b.������i�$s���!�e����k�ߒyew�@���s���' �iCa��$͖�_J���w��f-IW������&Bk3��f�g�KO��Z���Qu}zZ��sI���r?�9W�n��H�Y�A�#�\o�؅f��s;2�*���o��;��7��N@�D@gr`S���+~ Zh\\��סZ�p��Ju^�z��ˊ���i/�I��Ռ��F��@����2V��<
 ���d#z'3����>q@�i�'�����*�ŧ�[�AM���Dl7(�W _/*����&ο����S�V�\1����	�NMպ,�V�����t�`I�3|׎c����Oh���H���� 2V���,�zA��-x$7�1A�AC�:H�*��ǲ�Go�f�&X�T��Y3�E{����U0�>��.�l��M�9��*0��;%דL]���;Ui{b�,���Y�������:m�l
}l^ef�\6�9��*�o+�x;X�V^]/������9�h�}@����R�ю��i�|c�D�
g�+Ͷju[�Ρ�E$>�O^Ͱ�f��a�).�[���ť�+��Q�6�$*\��� ����e�	��y'� fm)08���A�6b�E��	&Q�������88A���(��C��O�v��[���j�zzi����E�jS-�dB+��xx]j�9�F; -H�S?���8�R�}�@���dL�QWl#�vv�#��^Npcz�j��ћ�8//p�,k�+5/ڒpYj~:!��ѹ��)n�i����YW��F�`sݻ��,O?�?Xt����+ϕ�m��_ЮIvJi�eZ�׹��I2�
0�Hv�eCѥ5x��!O�]cK�#�-qٰ�UCI�i%�JAtN-�V������T����v�X��F*[\��uI�Cc:�C�\��G�B��0��&��A����I�yH$�r�>�b�;����aK��,g����IH�4����<��-=��g[�K&qX�wK~�|$3о�E�<^Iiq{w$W��7$N<�Lι�0{��T��i�P��=�	eu:�.i�=�B;?��GL��F�fn�:�e�qM9��X�8'�_�1�j�� o��SFL�3������������s�q�2�agl���"��H���1}�->���>�A��6�
f�i�8��[Zi�F��0	���1��
���o�7i��-�㌼�|��#cyj=S4�½�Aqb��Ŭ�{���_'��|��mYa�m�WW͑���b�'>����yH�j�[��u�`���Ԗ�9�/�>lQW3mY�8����8���`���\��4�6'X�WX9G>ԡp�x���%6f׵	Ȩ���[qѡ��=!Ց�G�x��� ��>�:��˺�SU���Y�5[{�������T��uW�[��,���5���6�MD0�yn3j�z���ʋo��)X�g3k폪]U�(>6�#'A�|1Us���l�|� �%B�F?dT�$�CҾ��(���d܄Di㌏���Fx�q�Ë�J�81鶴����f�%4i-֪5>w&��`O��x3�B��ʧK\kjS�� ��429��Ċ��~���T˃:eT1���H��n��ꃩjO\9�l��b��㤏�iqR[c�=�wd�t�=��S:������mf{�1�(�;�@(ֆqp��&�5�V���ơG�]=E����[�릭�J�e��5Z?G���.|�e�����9Hѝ�9�I脖�؁���(��QQ[�U��w����]̽��=�ȡ�^W
G�(�����đJ�sb�Cw�S��m:�������7�1���b��{�܍ʀ��~-G�#��UJk�b�Ǡ�U7��Zdn:���[�`���swo��Y�R��pp�9l��� ��In����+�Q`m�$w�$��*	�a�E��u�M� Ƣ�������q�X��퍅�>���=��)g�_^�PvR��0z�<b��j�9TH��N���TV��p
��_��h�MB��!u�om���>T�M� ����uL�H�s>�sa��c!�ޚhP��k(`O�����^���Ԏ��t����HX��x"K�����^"ry�ǣ�S��+u���q��O�:�N�wG1+f	6�%8ɹ���L��_��M��W��{�c�(OD}Z��m�����������E,���A�J���㾃|���qJ�KBE�װ^�4���
a�+?����.��?���x2w�	O��vi��h�Ug�tWg��&T�H�d��4���h�}�لO�ϗE~8/(@�U��F��	*��.N{Yjw�k|���]�R��ܽ+��G����J��]�p}�������46�IY<w�\/o����_�O~v�^�RLz���8��nᯡ!˚[Y���3���Wo������y�X�I0�gd"���9�kI�K��p�l�)�����᜼~b���o���A\	nS
�4�i�-��ed�?J!+�d~+6 ��GbO���ͩ����nS���?5���	Zu^��T�D9j\��Ȅ��F��m�&��88'���� �j�+�
Dy"Yq�d�"�7�*���	XS��^2P�}Cr���	�<��P��fh�흵�X��O]�e���8�VsR�Ӵd�?�ջ�	����t$n�&\��G|�;�XY��g�V#i��##yz{/J�����&�<\�~dV�9E��Ǧ�=�vDgO�#l�j��C"f��>fV��0js�m�Z����`V�)�4NF�5C�my�Wqb:����8���Y����rEp4R9�}{j<��:f)�i��j	&�Z9�M��
�ٽ�}�h�&NT|gԂ8Ha�5�����t D�G׮�������e��x^UKK�u,צ�&7�a��=�P��`���b�o�	�yJ��ki��d|�X��K��?-U�Vtzx�JzEuW�Y�1��-�ԋ��_e���,�	�ך~��^߫z�#;�O ��Ϊ����<N��$!9���0�q��x�Y��<
,Y���u�i1���Y��m'����[L��w�u؝�Oɚ*�/I}qwlby6��~t��t�[���c���d�{�i��t��\ԯ�*0�ۢb�[O�/�;�4`[n�ן8gh�ǸU&�JF6��	���tL�Ҵ.�`!�U���tp&��DжJ����7k,��eAX��|'xNz�-�~�m:����^���Wz��d�C�ʛG5�8%�|{p��>���{�N.��a���M�z��A �y��(�]�7�$K��E��K�k����Qu��9|�E#QX3��ձ����U��k�`0��I\.o�O��\G�j��e�(� 5�����dEε)�޹�z_|:Spw�%I�b#��k���UTq�o9K^6Q�+��_�K�󻟸���BWQM�pR@%���\W+����ט��y���+-Z���y�Da�6���uBj�Th�Whes ��[�]��2���8������>ϼa����KTB�\�ќ�D��W��'E�G�z��G���E}�k���r�����_^%z��xy���./<��n��s���.zQ������%~Ȗ�RE7�Ͳ�a��V�
�*�Cy�0����OPNucIm���I/X�:C��3�4SQ�ot��1�!	�>Z�W-��	|�J��C�a�ɮe^X;1+���'RLoCg�=xz)t�"���6��H�l��+ӓ�KK;�^J829�������&�|�'Ͳ�	-�S����><���J���@t�T>�$n�x�^�VKhZ�&p܈��3�j�%��#*y�~�4���K{��'H�=�t� �h�B�;M����4�9�f����u߃�8�.�T��� D8+���ҩ��;5;f=	��.�%VW�%(�b<xɡ�\�������_�i��jp����Vi�*,�D�3ލ�@�uAR�SU{|k�V��Ԕ,}PZ�+m��Ǻ
�x-$�hj�� �PƟf�L��YjwY�r�h��c����;�Z�e:���g�d��E���Zz�Wn��C$�[E ; �u[��$M������e�S5T!*AB�~g>O#7��V��d���_�.�ȹ���<�m���`��o �����6�����2�*c�.��,a�y�B]ص_Y�F��3
����gu��	<�Lo�2�yu&�G�o�z���P[�W<w��9���M�}wH�uTa�!D(70������2q����]%�i�ll���<��
�p���|¾]�1�X�u�_���7o��|�R����.׏����R�;(��6Z��?���-&��!�hS���r#�h=66;F�05{?��:�P���(�KL1���X%��Y���`�j���s[���@�x*�-�^��2���s����yav��B%����x������R#�7�l<hg��tnyHlιV|܅V<z�m��U1������A�����Ze�!�L�s�)S�18=m:���Z\���^��+�}��Y����hH�>ˢy6��E�H���|�`�;�k�[/���P{r�ھ�=s������eu��Yu�7����|��"L��c	4N��uٹ�zḷ�A\$bT������H�L�	֩�m?:�{3ߍ����ax��I��hA��e�E�`�c1�9$���鏠ڼ|Xf�`�g`; �0�y����^���Y��_Zr��kFn�a�拘���ˆB���pCoDKe�l^l���+ߓ�,���2.��~B��x�I3����زe�d��:�k�{�t�6I4ㆽn6����Y�9���VU^�~\��L�O��>�`�!�>0�e�{�T!K�b�����v^/R��?�}�&��}F9M�:��ƭ-d8N�k.eºS!�u�W����RB��p�0���2�����w(f9Vbx�������!e��U��8�7���
ߜ�ä��kf�����vt���03��<~u>��r�I�����t��u��h���0A��(��o�Z��n���~#d�bo��� L+��>պ�%��F�,AQ����O�6����%Z���R�H�v�+T�b������yM[��$i�A�6��Pc�\	O�cD���jZ�����؇n�)Ga��D�a��.�邼�GMj����5�����/^���&l�7��M0�\�.wqs�m*����,(-%���b������Cr�j��P�p�5�4q"GG�������gM�0��y�*w�8��9 b)U�|��,単A�a�J+�G�춖�LX�xY���V��o2���������Z�|�v*���v?�:PGI��8�k�a���l��a�OmyY��?����|썢"Td/Ky�@���?Ϩ���S�]���2�X�]+1^O/h_���>H�� �n<�G���� ��'�0	��?)1��O�6�</W��w7��"����hCH
%;��U��TL3�P�2���Cp���9�P���dz8T��;q4џl̈������o�d��)j;O@����O5xL�x�T���u��p.|��������{�B�}�d�����ꧽ?kQ�o��kyx��vw�ӥ�*�:lB�U��Ѩ��|	4	��3�^,�s�#�H��3M��͗�8��֦�(@�{$��L���5LY�$�9��j�սhQa# ~��f^��@��߳��?�}�<f06�OzHsLz����Ķeg��Y�Hx�`_�'g��}�9�f�mߗ_�cQ�X��M2�#G�+�=+3��3&��v���y�h�9�2�����
b�� e �5ˤ��HC#d���HE��0�##*C�Q�ѷ��!�c>kS8\��/pd��o�#���r��?,��սh����7�i��6�y:�#�����1١d����ߞ�V<,{����n_�Nq���n�W~C*v�/��٘?�;��� W���0��{��)v�)D�ad[\*V�ǈ��Cx��Q��5;}ѳ�r�T�����,���_�9���y]�������A�zf.Jƍ$�LYb,ꆲ�L�j�X�i��/�4J�4�����z�Ѧ�݉'�_�W����ؾ#����npq��"�i�X��`UU�)e=�u4��J|y���;����l���Dɉ�H�?d�#�*���Q.+
X+!�ꥬ8r���������%m�H*��nhKӳCnA����)	eN����b}�3y�V���ɰ�"���!�֞�cj̄�By�w��A�m��l�57�\d����wK�\��w�-���ߖMFgѷ�Ὕͮ��%Ãx�o� �֓�}�e��x��;Oӝ���,�g,�$���S���_��r�K�3'���?G��_}�ok�z����
O�Z9��$��IDa-m�i۝-A���̬�����V�b���?.�<�cg��C�j�������m��h؆Wr���|��dI�{�����+i6n+�[	��0F��[+�<�s-$�iG�`-�qAm�]���&J��ȿ�>5b�@���6%:�̲�Q2��$�.��Pg�3Ќ�|�%X�m�'+|�m�w���u3�sʪE�Nн�/(��b�V,��%"=�b#�y��Da!�:ō��/�y�_h�D�6�\��3�cnJ�K��F��&�_��)+��F<��f��y��w����/X�_z,rYÈ��(ۃYk��V��(��>�r:�9�Ʉ������˺k�Rg��Ƞ��/u[7����ɓ�i�qڪ������K�pIV���:���h�u��;�W��:���%.J� ��\$����|���q�ъo�)�j����*:k�{�UP��F��eV�V�;O������@�~�j��u�?�+&j����/�2.�U����>e/�J4F'Hh������J/�ݔKrrP��_��M� ��W.�x(�XX�H�6*��A��.�B��
���^�ȓC���S�*��Ҳ�d>�Bǥ?yO7cC�d\��N�Wn-m�RuIϞ��H<����͐Oe䞚|0k��{ȼ��n�?��l��;��60���(�E��OtB�R�E���R�o��BBCaD4?��#���qg�����:P��_���jA0O�.���7<��d�1���@���v}}}�;hո�WX��^����xm՗�>w����l"�)�ܫ*��S�W�Z~�)��c�#��A���x����E����]���:n��̊D�+[���e�t����%�#����+�VO�H��7"�X���ġ�}����>���5�BB�u��t~/�k����e{O�����>�WȺ��8d�`Й�:Uͺ���ڇ ���-�?�J����L�gd���%�m�`ѥ�_J�J4��y�-Nʖ����#�u�{l���I3��jx"�9,�b���E�r0/V���`[W������� c�_{���f�ũf�L J� ��Ε�H0�,:��c1�@m�:"%d7���A��SgL���;���P�L���V��Z	l�k|����X���������T�
�M&��3��|��6�Vq�g k�P��s��ۙ���Ȁ!_?@5��Ϳ���@
�O�(��rbDw�j?�O��ex��B��e-�A��ALD�V5�[T������4=�Z��>o lD�;<�x�������7HW]H�^>Zѐ;��{e�Ϗ|�]��DC�=a�'T1:��#	:
���8�x~�9�]�����D ���4ڴS��&���ŏH@����-�
I>�įn�y���2�{4ɠ㵹�2[�R�{(�9����l7]�3�����z���?���������L�s�_U�Wxd�4�ql��;���ӱ���͂� ��zx��5N�1X?��kP��B;�N��h#�15��6A�k��zV0������Oqݰ�6L�e�At#7)�]�U�"Cօ��h�B	��_ޔ�W�r��'�����U��S,踻�P䵠��Hk�;�
���c>][1(ƻ�~_%�ZԄ��gnq$��y��9�$��J̖��F�#�����!���)ۓ)U�e��'C��c^�3��:|���]����2B�`��:�S�(��*z���ӻs��M�H�otm6 �K�8�)%���@�JFGw�	��p5�@�ǉ���Id)\6�
S2�������������I�
h㙞��K�7v�A*_*��t�ݩ�@`���*��ȦK�rp��p�I"�1+����?Xw>�3�Z�n�V�P1���gO��'~-�~����B�!n�K�Pb�k�ASkX��S}�s�j\���e��g�P��@���������m�� ��[��7�м��λ+�{�?,��� 삢��	(0�5Hiu�X�w�xK�s�GTc�'_�M��\\���u�7|�L܄#�t�0��Ӌ�>7�~�F��wr/3]2(�*a�n9�)�	�{w��L%�����L-,݂����%�%,��S�
�f����o>�7�>w
K���k�coMx��,8�"����k٦��4"�'���Z�?�}�sc@J��}�ӵ�޹�:v�T���C8;��DEᣱ7��Y� t�ĳ&��Z�,w:��;��)յLj=�Zo��f.y�.
��I;RCu�a���)���cA�u�ZD���]@��A��퓁l�u���R��~B�_s���i$�QfFo؏���_ME�I�>ˢ���GLA�NX�4jq?��c
#+����q�J��V�.,J�bX�"��y%���� �xT�7{kKB
2f���̅6��imIo��PO{q��ũ9<�	�Q�Ŵ �O��q�L;A�e�oh��%}��Z��pys��
��|��M�8k�Z��� ?+�_���k��|��÷Tg1�{YO��_�EwT�vr�BZ�(CA�T\����ne�RJ�����ΐ�#�]=�K�j.��m�n~�O����U���o��x�t���=
����K1W��ˎ�Hܬ����4)�U�����?㵯�J�)��%.F�:\�e��Tmq�L��/`�`�ձ,s_�_���	�6� �c�d���Y獢(VqSq���m�$���Ã��'�T�>��z-��'�&>`�X�}�b�ų�H�������w��	�]�
���:H;�nלQ/n?�l㾐��d��O�l�����-�'��H���`�2�&O����^�E@Y� ��!�?���%�v���c���a_cʼ�m�2?3@|Ց����	�{ֿ�0OEn�Py�����XLӼ����aUu]�(�����F��S����n����;	�i8�t����������1ǜk�������SD!߅�����#·mp�@rc'�����*�w�b��C��b��I����$\c�o�h2gN�%o՛ɰ�~��Lm+�r�<��b�/��؍s!~!憑���bg]{�8�ރ�|�m⽇�y~�ݳ�vʣ�S�O$�;��a%�Y�`0u����1��>b$��L8$H`�'0!�7v���Aէ��r\!Y�Z2�{��5�Jd;?U��4�bn%p0�4� �W�I#�F�Ӣ�(B���X�r��V�	'N��L�ע'�h�`��K���4�������kT�3Ű��x�����/<�����Hp�
,�FO,Sw��/���w�
?k�IV����BL����r���e�:A����;�K\�0�����a���?�*��<21� oxY����++^
���a�����6M�>uC��Dt���I#�A��&b�M68 2�J/���3jT���].E)�͉4o�cC���C"��`b���3d���k�%��\]O:���Y�5@=�Z�^py�����5p$�� �����Qy�?�z0f�7�����b�2�*XS_�p�e;K��H�b��"h��h��	
��f��x���,#A��ظ�q&���W6�?��[�P$oN����z��s���fl�<uTx��l?i�W��w���乭�X��GY���k���JR�)3����Q��S���uR���hQ$*3���؈(�d�>���lp�+	�,Tm��sK�CK���z�q�Q�ѝ&�|`.	������n�۴��#܆��dҞms�Q�Ѕ��X�8�n���M���}�u�1�:�~��6G<(<��B)H�3�5*(ksQqK�'����J-1@�t�;o��159�������-�����2���N	�S��$���}g��D�%�y�r��@���"->8���e�I%��@5�Wuq;4#~��	|����I��W!.��x����gW�E�����������ɸ0ZT��ONA?ǰ&1�h� Ѧ��uI��gHoG��V�ܚ�"��o��=�MRWIW0I�x��V��'�T�x>���Ä�{%"dN^��>J|�a�;����VԵ�:�i/����V�����y�z�V�<h��iƮa1_�~ɉ=R.�z���XQ9�k��͹�VX켓�w�������~`AL�*Q'�P������k1DH?��O��/]�H�8�kX["�=�;�����ͻaY,<x
�4�Fy4;�Zk�;�+!�r�� ��0'�p'���~|���/�������}�* ���1a5�*�ɦ��/�H��E�DQ��5g��\GuJ/�YwG��S�*N��٦�Pfէ0����t�(�Ǻ3�����BA�I��3e5��P�+;1����mND�BS� �I ę��|y��B����[�*��ɕ��p YJ�_Q��ۋ���?�+��w��^Tw�|bX���\��Hv�j��_�&�+*E(��m&�>[6I�$��]�(NnK$���D��C.�S�C���K)�X��Z��Z �I�W�(�bb�{ӏ:��zw0�Ҙ����YIOc��лW����c�8G��ۼ{����Dr��I���e0�y1����ԉ4h��fP<����I�O�} ��Ap	�}X��K�K��27Hz2���!�v��2	��.���$�Y�5�;es����Q�����,h{�7�*�A�q̷��ҙ�U��dT�p�:��$ÀֆLy��Ӎ�P�ͬȰk��%���a��?�fVɪ�Pe�,���%����3��l���<+�Ѳ!p�oh56�X��
�����i��G�OI%{*B�/�f�^�qd�w�EYj]^/��3����������)�i�%9�����ެ�b����=)V�f�m~���q\>��0v����Y���)~�I
�;6�����E&���ϐ,��W�4�/��y�̱�]��X�h�� ��Kc>%�R<`O�^���׌������1��w�*2�p/�-�RȂ��cͲy�z���AQ@�E_p8Ep���/{м'�T�Sӿ�~�hDPCbH���;g�?`�s{��Z���A�ѿb�RU=������J�O��i�� ��i���i��s#�=�������n+��J�b��EO� @c��髓��!Gs�04��Rj�GШ��wû�u����e��/+�& o��[Y��x��,�♛-����pvP�!?��2�QM�:B���Ârn3��|��B2�c��7� ��ݫ����p�n��^C����؋��G��y>͚NQ}S|����0�dTe��(6�L�?u��M��9���lE������Ӳ라��oE��!������ʢ����We�S)�p��GF/�+&̋�n�v�s֒����
�'#������1
T썑5��A�oGz��*B�*�>�K-�T0ڐS	
@_���$�S�ܶ��b-fr������i�+�/��� ���û��uH.�E�KP�"=s��`!�������
N8<Q�&��s�9����m��8��J��.��
�����j;
ze���gWU�<n���ִ0ە7��1A�Ր�#?+�}�l'�>�́�D¿x{�皛��ڗ�{+:"W���:��E�h���\�!n�||K_N|S!����� b�?���m(�]�~t��V�F\�IhJ��O����j�O�Q�[�0������=�[�EN���B
��U{�-���^�R#7�b�|J&��,��9ۘ����ͅ2=��4�ԯ�ԧ��gfB����ś�>d��0\#����{��A�ω����O>V*��K-\v���=�ш����Y���)=��?y!{ �Q!6&(����y<�CZ���'��y�hj"�Jl��A�&g���I��{���EU��=٧�ּ�\w���*/7M�Fϟt��΀8)����^���@�:�7�7�/1��h<�F�Pt:�b)i�1,����:�z�AE)�񺁅��%Q1��a|L2�D/�1�,j �Ԯ��� oY�Z�YHF6��E��R�ݜ]b c�\��G�����U�C����V��8,�)�1F
�s-J��5Iq�B��dUI�P��s�z����*�BAfoݧtj뗖��K'�����Zq�oIr�}K1�d�~�P��h1eIB��G���/	([��f~Ƭ�
� ���c��ɢ�
�����G����M��*��?N�۸�>�yr��ڑ\J=>_.�@��D�����$� �EUn5�:zE�0�p|A�'���PƜ��e%��'�G�E�<����sc^�ߋ�32���c�!��$bI�:���|����Y���ެ|�#�R(��B��J&m�yF�4W0
���;05���j�o`��p�ڪ��@�&��������t P8���QHd�Y���σNu]�b�j�����q`��O��oK�l�!�5�"t�G��e+�:����/��g��Z ��!@�ʑ|�(p.BOzZ��:����Gm�ɽ�J�sxM@����g�����ԓϐihI�2���p?�քK��7M�x ��ֻ�Ԡ�&�o�6��L�+Ƴ��P
��?-����$��gXv�E�-HP>����U�:��MJ�(}����WCV!n�Q�=X��6'<'��l�/*�[K�7�~	�ه�
?złP5Ӻ���f�}r:HKt��![���j���pO��I`M5�\ǋ7
�#_˲�r��n��ک��'�'up�>�����>��3|����#�o��D�Y���{� �k:�r��0�)���"�R����MU)��Jl��S��;��ioH�]?��KkW�r��}+�v�����ىT(ޅ�5�ʹ����"�Հ@R(��P hi���j[��#�7�0�c6�����\�hP���}1�J��sa�j@�eCz���x�Q�i����KNS��j�V�l��п��x ��[��I�/�	i��W�O$����~I���͊�O6࿂�k�j$��V�DãdJ �L���ý�yM�/Z�R[�Qٵ)gVQ�I���o4��88T��� �㫿!��>F�#7?S���4F+�#�<�M����ġ[�A��b�&@�@|�(��1��/3'�j���Z6����|��@�<�6�s�B�})Z�X��%�a���%���DR�!+�I��7b4�3�����az}��_@{.�s�ia�*�����qX������G��	 �&��/3� ����A��2AbW�s���-va,��c��N�׊&���;ai�^/'�Ǧ0��1d ��~)�#V�`���A���5���?d�[So6Kd�߁����^�'�9�&]w(o�%��xPL��RidF��u�)ѭE��l.�*�q�Mo�^G���Q�����
�Ь�{�ʀ�_�)�7����ķk��)���0U����
"u4�*�"���W��Nz�/eř��e�:�_6���ȩ,�ӎ\�~5�{$�����:�/�.�����[��f!uH������'{��Z��!�G<��
i�\?�P�v���> '�%��y�"�Ev������
� X�$lr?"��~�e�D��ȷ�"�k�_����,�uh#�>�N��@�������D-�z�Z��=�QQ�;���TzT��|�\�U$�G}��u?�[�L��0Ѽ�ǅI;Ev�TT�F�m3[B�v��Oe��e- 8J��=�D�~luԔ���Ǉ�I������}�ͽ:.)�Gm��?��I?(;���,}�	��}R�jY� 6��� bXb\�j�A������-ژ� ��O@�&��<�#8X[��Gz
��Eg>�n��V�\`��/<b+�E*6陆w�#|��o@��[t���M�*�0rc�5uV�����W:S��	���~��+��X��K�� F49�:�T|^_�[((�;�EI���p��H�����ݯv�J���!sh�N���%L'ʅ�h�\�\��/J�(r�מe�h}�EӨ)mX�Z��U�wU�&�o��P��
�`']�W=� .L���&׊�o'v3I�Y/7�!!��D�2h0�Ģ`�	�.k�R�Fґ������>=�������K��U�6cA���ׇ)|P7�e�3,�������ҤJDザ���\��-ՠwV~����P��Nu	/#IR�.� � 7R��$�����!��K���$.��X��Oa�X����Q��k�����<ilU�l������+�Z�!�EP�&�*,`*�Ͱ71�4oy7���Y<���-Ʊ+�6�j���b_,�E,G>8��Paa��S}���Z��B�7� J���Ux��MU��������>��� }M�V��D�ֿ9_{q_H����J$������d�S ]�Pa�l������
|x�Tp�=>[��ӭ3 rI{T�5����O4�s�P��:w��f!�a�8�A!v��}9���*j�{��խs��*�\��A�^V��TG����G�'/�􅘃ฏ�����12]H�=0]Ki~ǿ����z�/iK-�����Ađ\s����=��e�s�����z{�ˠ�>���b�w��������Fx��� ��&�
�N�'��a)\��Ϸ06�(����-6_࡝��j�?��@b�J�,ׁ?��r�AL��u�;@�t��/*O�R�p�Cw�!��4.�z�m�oH�W��ST�Fo�XMi���5N��l:�>♭�7I�
(�$�����> 6�/ M�W�x���o�R��8��9)��A�P�uY�5R��xeZc��N0��_�g�B�#ߩ��$5��\oR�M���X�]����8П������TRl^os�,BL�}�q��Ⱦ��T~"���᫠W�+��6����I���)�N� S�]�a�;��$���^��} �T�9ej�>b ^b��Z���v���|��$�}��ΣCc�Sm�#��~�Y�V��_f{�z�
����F0���}�:���i�ˏ�Oʱ�,������^��D����0��� �Ȳ/�|��:M���nn���v�P�M>a����\v�5_��6x<h�@;���PfI�-������l�^�=B�{{�6� ~���I�!5���:I,-����
�����kAД�J�(�x�JN��/�W�-+�A�ݽ$E��l`
F���	�\���9������o|n++����YK-��L;����E�]?����c+�_cYjb��/bG5ZY�%f�P�F�&|6|Q.���y�`��ȭ�C�wU�thxYS��Z�u���b������
����^ap��H��J��9���`H/p��獏G.:�헳
b�N|@y͡�@�~�X�z�֔ u�G�B#v�0��oz^�wR6��/�����v��t:��f,:X}|�r�w\���!|��� *3{gl)�z�!S��YH��W�ȶS�fPBg+v���"�!2���M�F'2�!0% ��Yuɯ�{���ݽO����b,oa���D��^�(�|��J��k�K���)^׃�OWQ'ӵ���̷�c�
�B���OE��旒���_����<Zɚ�D�v�evά�
���<�c�(�h��gYzĕ�2j`Sx��#�����U��������u0jD��.8�+�����l�u�+�@���{�k��[�G
������v�Ů��Ey��<P.Z$�B]��
����r���x[Zj^8a�������oe5���,yޖ/�`.e�ozH)k�'�+�B-&���1��=#�@�.��b��JT/ɰ5J�;��2��]�>�ca*� F�w��t�\(q�%U�.UYZ�U��2�n�Y����u$3}v���2]�SWQuJ����]a��*%�$�g��]��H�l8[��w�w��H]�i��Wi`<pf��~�	OYjl���������l+�a"�n\�^Y/6�}}C�}�H
w��lV(��ɗ_�6��M�sr[��~T�K����2�����D��R���_��D?�"`@ G���(�pɂ��ۼ5����-�x�꿨{�	�Dk��;��Ex��R�צ�Q�\�=�V6ʢ���|��P��gd�(R�x����u�����X�w��v^p��Y��>c��s�NG?��H��ʊm�p�YP�H��N|P@��o?9Į�ƸϨK�Ş� +�,�d�=4�n=P��L�dQ%~�}��|�I6z~gUu��p����z)Wo��I&Ŗ�Bs�W�⟑�GW���p>�ڙ�b��z��b9I��D�45�&JB�����h��2A�[`+3�@��B l�7���"Y_to�ϙ<s�$����b
r{=��[ȌѬ�4��9�ù�=8<�;�8M�ݲ��;�ؓ�ǹ�o��Gb��|����֏���C��������@�?�U��N\��]lE`����E]u��R�L�/*�T|�_1fG}�c��,u`|~���<o���ܬU$+�?[���zb��k��m��q:yݷ+��J6�!ȗ�3�
Ė���"Xj�y[ ��s������~������`&DP��ޛM���s����*N�퉗U-�X�]�P,��y}�����g�2�$�tqoV��ǿ,u�[fH�/��Nu2AZT�%tH���>y�J�ց�x���3�2���g���2E Ěpz{/'�:؇׬3���f=3aBG��Gzu�cC�����wg9��;m�-4�(i�����P.4���wѾaZ1���@�w��W��Qi�,�K��H�~՟Kc�!�iM��%��L��HX��p��fT��B�$;�h�!���\K0�{`�\�uۓ��l���J&������������N�J:Y��01��J�l;+�9l�Mx�:S���r^�PB�?(�D��
���R���!⾫��ܜ-�_e+�z��W_r��t'�Ih������q���Bڮ-� ������{�x:j��a^�E�(����MQ9���Rl��#��%�RlƄ��$�B&i�b��ߎ����]��3����>�WJ-��>�֛ܽ��s�����&�9dJ)�ة5˲�-,d`EUr�еC�����GQ{���?�T��%�g ���Ho��b��wn�+[l��2���Ҝ��ϗFp������8l��&�.,:�����!%ߙ�L��RC�<pa4��; gW럾Jn.���uWq�5�T���r�h�>�p�*��9%f&����|���M��XZr��jzB�['��B�c}�ň�j���.�j.�\+6,,bb���#g�7����z�	���7ci@˯B�:�`���B%�#����l,=&h��n�mCף��M��t�n�xh�� ��L���0�	��~>���F�W܊��Vf�T#)� �԰�b'wz��U
󇶯a}����^J�/�[$���������K$��|�l6�u3��w��.Kh�|4̵�� խ�4�����Vk����c19w��NdzJգ��3�2ת��q9�����>��	�V���OEo>Dƈ�!�������֜1J�a#����p�{�^��0��qr����0��p��,�łH�~����r�81q��n%^]�!j�v�v%f16(�V�{��D�k\n��r��*��n3�C��y�X�!�`�͵g:�>��B�a_6��К"%@�Eitم�n�e�u��������yb��F�K*�ԭN��p��� �"������۲�
|�+��ޢW�:_XC=��E��uj7�~�ח��J-f˚Q�j�H��k��z	�İ6���N(õ����4d#����q/$7P[3;��I�o��W��Hj�#QOS��`�N�\k��J̀�_������߅�%���,IM��dHd��@���C�M|�ˀ}�WS�;�|^���`�U���g�|�/���mw;�+$n͎#8'�x�f�0&���1B;c��Q/���R��M�KǴ]��]���o�:`�f��A䷠���.�������g���f}y:U��t����m�Mq������Q��,�g�E����eƈP'��Z���H�`'�C�c����7s�%���4�VzX1[�`ڋ�cI��#�L�$��t5&~u��'��%O�~�g,m���x���b2���]��3,�d�Y5[her��]�ƄZ�A�����w%�����\̝Tև����_4)���4�7��!$y���1�:հ�����e8y̵�y���Դc�{خOS�l��m��@�Z�qHY/P!�s/�10���R-j5��	sLx1�?���e�C���K�B\`��܃~���K}���^C�9���]�)�t���1�j*�$�IlBɡ��!��y���L��qc��I�a��~�>��6H��L���`m���Z9�?2�x���i��w����5��i��ĵ�v�l�a�>��3�EW����>�}l�v��j�*���C�V�
�;���ٰ墼 (�cm61�H���㘙g��*�<��y2q�O�aŒG������`�RY���i{m��}�y�Ș��x��O�+��g��SJ=w��'��(|M^��*�H�.���wK>�!]�t��lϬq�81�������Z��D��&+��*�^C��N���U3r�H���w�4�ڼo�#'�����Z�M9.�m����f
�)m6'et��GL5&�k��,�T�^w�S���4�N���N���!|�2F�=�xܗ�8(6%t��V��N C���Ah�� u9���~��y�C�4n�������v�c�٣��MG���oG��`Kߙ�P�YgH�|���W��W��ƀv��^tækq1��Sjn���5dp�敶�͙.���w(��"�ίF}I��Z��T��h(^K�E2=qX��'畞�\R�	� l���Sz(�n���a�,3i&yc�/gg�����H��� J�л���՜��-��QC�)^���yuoo=ws�5zB8y�s�ī����*�#l���Ͽn�1o����<�#�f�$�Q�HXg\��1��9>��g���\]���h�9j�j��1���"�|Ox
�^�N`�S�t]�F �C�_�c�d���o�\���W}��AÙB&t�]�*iq4����:���>���?����#W��k�Z�`�V�.̯�*�]
L�a�mM�-�k��NB����i)��e����U5�~;,��;̯�J�U�quUD��:���
ϣ|[���}��ɠ؂H gy��\*�LH>KL'Jj��"06�t�-+Q[����NQ���Ws�n>^FȎ�]�P���d_ȸ��gm�o"�HX�7�g�wg���q��}>[���p�:_V/4��f������6	�ġ��Be^Odp���s�W6����2�%���$��Nm������-�*�ԲN�Qp�����'	o�9��aR�����/*b��V�2�.��%k���y��$+^�r�݃�6�c��r��R�}����9���$f�d�]ʻ2�����і��,-e[����ɼS��Pfѻ��-�;��o���k���O��C�+x�j�ω�[���J6�W���t�{�͍���(���!�_#��SkJ�E�_t�Yh'��>�D_i�����5��M���@�8������_eO�m�H@��od��=����RԎ�+,�r���g���@�wJ���U�`�/z������=�{���4;n�����WN|��J��*a�_�ƒ���n���� fR�Z����Y��}���ߜ*#N=�^���:�Be�w�(�9��� J��,��Z��Y8J��<�\W�\xh�p��,��.=�&6�L4<�7����
j`ɬ�ݍ���b�lf����F�q�Md>�����0�
����7�֖��0�֕C�����$'3��f*��Ӷd�u��⋑E�3�e��X����&�z���I}���[�5>�Si���!�
1�r�UDC �! ��O�;���b�[��rڑ��Ά����#۸P� ���c[� ,�x���Ē�Y�/�^�`���Z8�c��_]!W�;�0 M{�~׉��4Ο�Q4�Qf3u6�k�����	. ���8ٽ��jOu`;r8YE��D��Z:1zU{�	S�a&G0�����AX���s�ʺ4��(K+��Iǡ��u���;��m���;G����qd���V��0���3�a)��]@���b�	K�p��5�ٝ�I�.���-��ҷ\-,�8��D�R�Q7�����q0��s��r):�L]\L��vey���DFG�N�Vv]uZ�߱��$�^	����^G���z�a驠tV/��a�/����q�������1 �1�2�6�=/>�m>�O�z"��%�f�7k�H]�oB^��0Q2Ƹ)�7�,Q��X��G]c=Z_�7h��$E7���#��$8#�x�~�:�8�3R~���M�>��ӈr�K�8V�����6:m�p-r̘>_s����{�e�@��h�����>a�8���MF�u��/&	�������dR���G��a;I�ل�V��춣��n9�+N��"ˑ	E��g���>}sR�����u��k��M��#��:u��axƂxt�_�-�dp����w]��uH�S�^u�+�@�:���(�vwʬ�E��c�~��V9%iy��:CAe�*���:Aam�agq�&�/J٦F2V��"��2��l��ڳx�/W����H�w��n����W���3����hr����j|�j�_xlz?!f�@�D��h�2p�\;V�G2�
}B�a�Ӽ�\�2���N<OITs�"�FU�L���yq��a�:���VO��a�ol��vJ)Z��e��`i�����Ze�{h{/1^�����F�Ϧ�Z�S���kH�A�)���B[15u���S�;ݞ�*~[(m1��-F0]� �i<���>p����Ԍ~�&��?�����]�x�Tt|8n�eZΒP���h�;��Q����8�&��wEM��`#1t-S�e�)�9���{�����
_�gI�̰���cx��K�1���]D<U�XS|�/�ғ)�%/�q��&��@�,�?��w�E�I��͙t��XL�����V��沒l�s	���P��α�������3���nS��\cq�|�m�������dZ�ǭ.����r�j��rkY{-ɜ�r�Z�,N�L	��� �Q�E�A���HFVieX�M��9�^F�M��U���D��2駪C�;���{T��ϔ&My��Qޥ��\�74k���h�}Zqay�?��;���T7��qz�ׅә;�����
�'Xn'[Rj�z~���,�l\gsãaK����	%�z��t1���I�C0y��.jϸ8�
"���M-R�ù���U��#����yg�I��s_�_x���Y��|�pF�CKk�S]�� ���i��(�J��W� ��aXb��z������s�|f=��)^���,��*��Ɗ��ڵ���!F8ʴtb����C�-��\��H]��~���@��A��č>�i;?Ō|c�\\��CbM��������EZ]2�֧����>;\�h쌗�ґ���e�<��������u�_�~H�8��Y�^l�I���j���D�^(3#g���(��/y�nscHl�J+��Oy0P��/�ˍ�θ�Ԥ���:'>Fx.#|&< n/�����9��aV�X��X�?i�H�*�m�!���»,3�1P!(�Zq$�p҆�0����n�)�^�-����[����CJ�IrT� ʳ����r-�U��CCT��0�Eq���Y�ow� .]A5k�|���>xC�׎UX�$Ԝ�Ր�b����"q�3�� �,���k8�w�-E�Ϲ���&����j�	|��v�H��� F�/��9k�'T5:��K�f��ēb��F���=.�Ն&���:�Os��u��AG	��Ɏ�۱�L4_��&İ���f.[Pj��6 �T=pXI�E�'�,g屫�V��vL*/N�D:���Y�1Y�g�8�����7І��[b���#J�a����l��$�oX��
�(��<d>g ����׉�� K�U,-��{�r�Ey�!z�A����,p���ǹ*��w��$?س����y����b����X��-���L��=b��Z�q�yx�w���B��U��&�߮�
Q�[�J�f���?�j�q;��qzw��9�\�a�����,�Ot!X
T���Z���� "2�ea'�Z;�3O���ϹB�}���Qh��u�1�c�<��f`1���9Cv���[���w��<zKo�"����ԧ�ex�i�ɹ��y˥Hh3+��8䷣��'�B�?y������pT��W	}�Ņ��beq�N��M�%��b;��� �� J�UDr�!&��GD�>Fd�JW�M��d��_��o6Ȭk5t[a�[~M�h��
�6}qDc���I�����/���Up�10�z3��&�o
v���+����-����� \�>D���p!9?���-vX̡u�� �SIp��������ٰ�5m��E�a��e����c��П��CVJ�b[.W�<���vϑߨ�Xv�{j8��,ֵ����N0��l㔶%�xM��;M��i���*�r۽w����m_Mf��c�l�%�+z���pa���M��w��Lo̿L-s_�{{⃿�����w5m����V������cП<u�UiÆ���>�iQ��
���g$MQ�X\$�R߹��BV��=*h	���<y�����c�k�_X�]���&@0������)�����;c1=�3��@�]�eg�Pxe�������ӟ���
|:����;�qN<���"Z�=��1������W�$m�I)�1���H�O P�|�jY����08�~:$i�I��<F7GOp�k����SĄ��6[� Y��Q�A��Y��`��K�����A*���W\c-�Ӥ��ӹ�У�`��˛�k�ͧTsU�NYz�\8Og�v$|ל�'4;��<)N����H09D���j
�8�eԵDG!��}�=��7�e���<sK6G�0�qbM��U�4��w�V�յg�A]�\��?����Ǿ�؟ $q��D��`��-���zcl�i�HN����.x�T�QC��+�qi�dތ֚�W#cb^����cBg�u@�P�w��հ�:��KQ7����sw����2�������Y}�E��`�o���zv�`�Cc����m��Q�۬8NQ���c5e������I�0-.�dV���xp*�h��p��I�Z���-�BfT%�_��8��R��{F]��k�������e< :�+�8*P�=f�J̋�����ƴ ����<j.ο6?���"��l���Y��l�}T��_�)m�>g��,��G�h��5I�5�sx��0���N����F����Z%,���J�cp[��)��RWT!�x�*|��K	/_� a��j�W_��C�dB�V�w�z�ֹ�	�S7�m�>�������FKZ�C�%�az^w���Q��2�̣����k^a���]B$��b�z�m[�4J/��^~ʈ���XI:7�v��C���5��6L�S��*Nc(��U�� �(+@$b�s{u(G6��׫s]9���q���Hs�G����O{󪫹�����hɢ+OZ�e}Ø]��Y�+�>r�9�w�0�N��AyN!q�MD%k�έ�F��O~L�u��h�d�b��]���1�X��Ӂ���t���p�%'L�7���8X�v�J�Eશd�sK�g*�ȩ�y�vd�>��zn��j���Io��zb �0�ۻ�R����l|��臠S�;8�N�2�}�#g��ѷ���5%�����#���À�m���Op�\��*4�7%2���ҡT(�|$�����I\{�$�i��׼Pώ�|��-d���_�r�����
D�W�OB��z���k�7���<�qL3�(��}`+ �+�&�������X���94���G}D/�h�j'o��{���w`5�z������di���"(.]yN]�l0ϗ!rJ���%�xH�O�t�9.��\Dkws�_��}�?�XXS��4���I�b#+Th}M�[�	���N���t�A��7΍�c[�9����i����K霼oh�*�j޲�\]"�aG"��"E�cr��L���b+K+�00E8v� ����!d��g�;f�ɆxK�?�(^]��;:���?�����6�5[r}1�a��h�YK�;n2GA[�ڤ�(���5�Pb�oq��s8�I�&˼��C*Z���_�8�JuC��<Lu:	��O8Cʔ����¸eX��ٜ�,������׬l$�B@��VA�u#�f������uX�_��\�~"��ߌ3*�z~v�<�Oȩ�.+��j�1d��12:�>�5]//�������O�l��h������Sⳙ E��r����֯H���[�r��Ǐ ������`"�������>>�Eچ9�D
+�5ܦ�I��J�ًi��j
�?U��!��ҕ{�Ѿ/-���eؠ1q�M�������Ӧ92SP��4ױ�=4n�T��ē�=�iE�J��ƺ�	��G�	�� ,+��77f�h��W��$&;ЉϡQs�f��\x#��p�O���0�������':*BFDA�(�N�M���BOX�pc���D;��yG4iR_Bw5]��z�2��J� Nm$j�
֑�x'�ţ��;����hc����Hڍ�]p�!y��h�S� �^f��\��͘z�;�s�tn9&����3yN�ҫԯ�\i�0�����C�ˍ=b�0nf���b�� �ax��� M��&�{��0�����鵐���G\��M�� ��}�A���E��UO��Z1����7cl�nO�`f�H6����k��Z��[�l5��&}F�
m>��>*�|�z3��n�'�YӜj���Ʒ�Н]kz�\Q��|x+,]��*�F8�����>F)i��:�s��b{ڛ�c@��b��u]�0�d\��g#/"P�4P&��`9���C�_t�Kdl$c�'7���"��3V%Y�r�����eG���}��֪v��Gԕ�����-ֲc���Z��U�aEn@�
-hQ9������	�;<��3c�f}��0�L����9Vr��Hi�wKuYܲ��k��؁ �F�9���k�Yn|�Ϫq��?�M���8x2l�Sy��a+��t�L�F����]��o�X�k�̐��!��jx�X�;�I��v����x�1�����k�#�d"�^J�7��*/�S{��	����&�a�pڋUқ��n�+q$�QG���(�H?eͣ���P/�Ru˾��������'�:(�vd�܂C$���?O	��������ak�$U��t2�ED2�A<��P1^� Q����֢^��!z�Y 0���`G��,��y���n(�JL,Py��m��|$�'�ՙ��c�8b./�j� ��s���.�巗���ǫ�L@��@&�O�<��h�5 ���NMd�E�� ie��~��Jw�.�I`[��,�M0�	����MW?2W��W��4��Ľ���ݵ�����+">�����g��*�4�<)�/�4��qP8�6�'��Tq!4F��
��U�Ɠ%|��!Rn�(��(�)�9���A�K��F�w�oN����qě�6��5B[
��9K���]�qH����
L˗����w&!��C�Ct��	f�EB��N�=Yd[b2Fy^�S��yު��G"��Ȏ����9aW(#�y��A�J��;�f�B��k��ڞ3��.j���e=XӋlIÈ7�f��5�|�]v
.]��G�WF���B��N!8�`�������������݃��vp�7��޷���Z�>=�U��vu�L����~��Z�JdXv'vi�a�]v�¶z�<����ɫ�(�$�P:���@���if:��ҙ�0��)]+�H���԰wF�����q`�]Wr���4{X��6� �z$�~��j�4�S�5�(B�Z��Z¯�r�ގX|�+-��"�j׳
 Pn���ϧ�5e�b4���.6�O��@��pw���F�{��{f����1��u�	��Eh�OWD�S���³�)����.=�0��~
,�(���P^�󂎰;5Խ�)	/Vc�>�������,`:����P�\2)p�F�~�u��z����
t����,'!���͵�Z����C��$�$��Q"�������h���\�tYًEz3^)�@aϥ��"�ԚmZ�I����ōz=��cg����"K/r%:A�5�p�w�M���1q+g� {�bҍ@8ԹO0%�fڙ���A�8W�p�g�)ƛ��j���'�_�EKE�Wi�A�K��"f*�{CA�\�wr 
�r��C��Le�M;M�?��Dߴ�Z=��{x[<�깳h�_J��z>����w�j�N#�����Wԫ���~�c�Mcz�ꪍ�-� r�Q[��g�5��*�v��'۱Z�� eDr�57�O���V�/K��:RK�O�V�7�W��!Z�
�OI��Z6�OU޷uK+������M�a[XЪ���vS, �;4�����Hm�pr�q]iS�y�M�����7�����A)���L9�ob����4��簄#���X?�n�\#��˯N��\VվF^T�!��77�?'k�LE���QA�p�,y��)���턄%�wXo�O�f���DP���"CcZ���0ts�Vr���}i�e��L7�C����w#<=��#�y=<A-
qOw�:�U�|c$��}�6t*:a���A��l�2��ی(����+�ց���3��Ӳ� $\��EQ�(g�*��+&]ƨB+:�f��z�
�xzV��A��<���2�/JG&���ٌD�<��M�&���2�"�ߊ��4�(O�)C�n�
a������#Y��	�A�Z��� +�Lk0��y� ��|Hn�N��^|������FE�(��T=��^���ằ��G �B���}��s[��^D����ݛ=��a�c1�5D�ޝ��uU����c�5��S����X͋��Ó ^�i��6,�%�W��o�ڽ
-�|G�C���H#��Ʌ���H�+��g�`����Ƹ�7�y�6���j&�}�P~8����aE�/���|3����6�$��bW��,�'t�!@�jb�qU�w��{ǹ N��b3"�/�K��㮷�υ�f��O^2�`��H�E�<GX��znѤ��v|s��d3��N!v�HH��2�͟s��p�2�a�����o�tb��	�\�t`�K�s�A���9riWu��Z�*�B�O�:`as������Zk��!��i�>��Lg�� +���[
�a1��
�7�ِ�haQE���H�p�S|��S:h�Y��_ y���C�o��Y:��+�1,��((�g������p�";䓃�G-7��t����;2�3�9�3MM�S7������}(�I�rV\\���$���j�_ތ��z�;q[�
�������n�95L�T�G��fd)�j^���&��B����DΗp=�x��>���N���q��<Ͽe��ͥ��މ��"�N� D�\�K7G���9���$���&�_�	 <��]�ş�����/ʓU���@��/]~sρ9��>�yA�lv�v]lB�<�;[����L�<���f,��d���X��wa$G%Lfٱҏ���(R��.A6�V�{��B�ǪA��ښe��@�Ͳ6m���?䴫��7�PR),.k���`i'l�ѯI&�G���S0�\xV�L�}�����@�]n�5�֊��d�������m.�[��?���������Cv]閠�:r��0�����[�b��<��U�H�*1�`�\�7��ZzvW�2�0.uHi�� g�vm���[��7�<��.��끢~Ø%Mg���D��\��y��p7��3�OY�K�a�.Mȟ�t<���Cq�.��/�+N׈�77}��?�1���Tp]��*!�F����Q�y� A��G[��Ub��Ɵgs���a�h�q��h�X�`7ۨ��{�]T�I�\��!F���H���H��E�z�:r�[*��i*C��vtFyz��#ukc?���>�ɗi��_�;��#�IF��B�4͇��fw��|׎�
�B�#��]�	�g�E�f���!"y2{��|�������@ �Pf7�������]�nb��0�s��_��=�*�m�W^��L�n��v���A��8/��ȷ� E�0��;��-��	����M��q�ժ�c~�9�����b+�!G$������ 5ryʧʪl���wE�3$�y=���ԉ�a^ĳ����/ՙO��Kr��z|���W��I�@9��k� (�̖Ki�T�2�}��hC�W�R�����t��N�����
��@4�vo��t��3}"����Je�Ϊ�Tи64��P���'٪G��߫�YY��>nWB�hٍ;�U�>��� �'f�F�Xc4��6C�g�Ӷj,�1�X@�e�n��q ���D�eOr��mG.��Ì�/����g>������#��L���a	�8\���T�&�<�	�׶Q��yC��c�}�ס���1����;U���S�~��*�<|�U|��գ���P�K���㮒��9w�΋Ȋ+�_*k�IK���+���꽘�Z.ܐ�������;��N�R�?��R��y��hA�\����=5�ރ��[?x�]T�0�Y��#�[�93��a����/S�@b6n��.*�<PǴ���*��kX/}��jM�C�m�����q+<���]@AG ��Ҕ����|uiʟ�Z�v��˴c�}��㗸���I�����ZY��}�H��-Г֞4ەZ��-$��8Ek�z��I���EBq������c��
Z�Y�h²�V�O'�/�(#�P��g�f!��&J��K�6�q_1�y���!�'�¤qze����3P��(̽�`g�ۭuD}����g-tZ�Fl$u��.�`�co�󾍺�F]�7��kئm'��am9y�#�r<c�*�������'�Y���I�3
?�Y�R��x	����^�����g[�-z4u0����<p�F���L�3r��ڲi��|���u�!�m�[��p&o����$�%a,��hi5qᭈ�%�r=�0���'
���=Y�-���B���qߋ=Ms����s;�:���16���l���/DAl��@ô�:(�@mV���,�u������T��B7�(~��:TW���r�;�Y�R&m��z��}kŷ��Ø�w:�c�������eQyh�A{�lV�h&?_�z} ���7�]\x�J�{S�M�#b�-XÌ���W��;|�� ��AN�����`Y������/N�y_>�a{�e�;yq���Oz���QX�i�{��ƥ�ꓞsrMUmť��D�qz���o��m��|�D��"��+J��(�/�V�F1.SF�U�$� �m���.�Ưb���~��WR^߸��qQ�p\P��I�����{���,)�7Ϳж�\��ݞp�e��U���^a@gf�δ+��Le�����:va��l(?�$	� ֆ�fHk�l�nl�v�e��\��k�y.a��I��4�gY����tC��kҢU�eh�ǆ��[;��{~�<cW^�e����L�Mc�Y��#}ՅUr��f�Tߩ%&��������T���@������p����WDnc�P@PV�Ҳu��m�}l�-��Q���ޅA	v�O�4� g�@�<b({-C}N]� O~qV���c�!������ɅB�U��������C	l��#�32,��g��c���#�!�4�$� �F�(Z��yHY�@�Dr�kC�T�
*+s��:��S�����!g5��R���t?Ժ�.�D!�Bx��I����o:���\wD�EB��mߎeFvV�s=���B��/2��P}����D.��Gl�ۣuk��p�"����3G5H����op]�SY
k����;43���q��(O8n���t�r��5�Wswb��ZA��[�Q*v*5f���"�x�G�j���E��K^
���h�4�+u۶>q#��^y��z�T%�v"�k��@�{h�q�Jʹr2�J���/#
�GZv�^��B�K��p�}�AK�0/[=w-���"+���R<��d�-O�_|A����-�z�%,�=<�8�ȮU���"]�������Q��U�nq�A}����Ƹ���]�����0쨷%�A���e�;�^�d���j���,s۱�9��TG��mZ���8iDc�� ���:<՛�>���YGmr��h��_���
n��2�>M��y�~�������}��|���?�8���, �����y[w��)=�����͵[�t�a�}��2_{�o��6 �<�#�j�eh�D�\?h��m42m���ݚ�8��������iNV���F]ʹ6|��u�Kj}t߸U�i�q�Y�T]?掾�d:iX��F~��^�LBn4d��8�N�^�l;��,����9��lYz�r����ɏ�߽��q�XG.m��&K��*�e���E��|�?(�s�W�b����`a�K(��-����{��x���
#�+B���_u7�،����؅a\\�$��"�ۦ�±e-�ʺ���RkP�y"��d����u���lB�_���	B����q�H���<��O����M��%��4G�N{�6]����wEUК$�2ewhY�sB6�������[0�X yL�,#;s!]���N�B�v\��b�>����H�$Sx;����ؔ�f�o��)����b��>
��bC�8��n�
�
�"�5����uW�J�I�\�߿�>掘�AmG	pa5͵S
"�DR�%_��gI¿j��0{N�Y}~�Ы��x7���w]�I�/��o��\[tfØ���0�l���]�7y��W�x��-���6�DM;���B KL�����Z�^_�x�O�$׌�|����!�sG��`I����7�V��K�@����e�j����g|�p�3v��QAK��$�ߩ�S��]�:���.�R4�O^jOj:=z�d�`ﴪ�԰vvu&d�i;��o���՟D��Z޹�{xF��Za��}w����{��a��Ϩ2B:���ۯ,4C��k�l_�ZRBEOd�x��3<��P�8`��V{{JwY��{�I<C8����Ƥ>Qx��1����2�W�?_>���M�թ�~�7�e���yy���ܜ�m�����Yu�n}���3e�x�/�c�QY-��(�f���"�l���ͫ"L�n�^�?��"x^α��Mٺ�K
ҎN��Ę��9q��S��*-ui���m�~�[<���#�L\�<��� ���y�E:5���%�QN9��x���lA|V�)�GX`��N�7��<����AY���1���#Ȕg+A��ʟ�?�x7{]�P�K��j9�pY��O����i^�݋5}H~W�� ��-�h�<��o���/?M��[�f#�5s�D �ۧ�v��B仌8ά>����2:�j{��0�Г��a'����"(�Tgp��W� :�-���D����-Wp��Sg@��K �\\*!�
�2.@v6?K.5��ז~�+�K ,���mxub�Ϟ�;�y1
?R�u0�ܻ��Z�,���ڥ�zͺ��P�F..�zx��i��x�R��ê����9$g��Yjی�=�����v1u��#�����#��Z�����J�w5۝�=P	��=�B��e�?�$��vֽV�i�K-���G�$�p}�h�Sq�{��Zh��GI��*�0��#��#Kq�����~C3�C�A�(n�[&�(������3�)��_�G��<Oc�i\^����x-Y�sB�S�����Z�ɰ�4W�C>M�f����R������+���շB���@��V��H!hܺ!�����W�o�k}>8��-�;]mٷ��=�y[8[�r-�����,֚n��O#	� ��h{�p�f�?ܿ}����z©>����`"8��6�K؁�G�Ϋ!�9227���ݚ��2G���zͺW�=��[/񮗌�U�d|;Y,+5�%�`�Y>�������RD$+�S4s[�@���J��b�s'�\s�,�M>���µ�l��v�-6;��E�o*����z!�L@%*DW��G��hY�|1"n���Ȃ�i�W ��D���w�"̩�@M��,�.m�O���$+�D,Orx�Xwry�w��,�����5H�H��r��Fx���+a?�Z;�l���/((я�Ec���z�U,�;Z��xz<�(�ڶ�u�6��}���%�r�	��'�kx�օ6�4�.����4"0���K�^�7�:�V�` q����_w��÷�+0�w�ni"���-1_�ȕ��q��;#K{[mfa��:�}�7��э�M�V;v�<7���ڊiw|M�����~��Y������u�;�QKT.��k�����?^]�S�
bC��_fv�)�:of���t�O���</;�������>����/9m���.)��9{s�y�=I #WD׺>���t��a���  �д!��Ч�)_)�aB��~_Fj̴�ڊ����1��S3������kc;VKE8������l2ԗ���^kC�Hj�˕e\p�'}~*���fk��#w<��)k�^�:�~��鍘��?|�jz��+(���^�� {�6��4�|����'֛�Xo�UVq�WjGcW�g`*���_F��\�E��M��@��m��"l��3������]ܥq<��>TW�[���6���A �m&�����^n>��Ƨw��,}��Z����G�����FA��7*�Ɋ�f�
�>|Z� ��v���߹����IR�7T(����������ε��(2�y)���2�w��XO���hC71�4�7�%hƸ,�=�J�iƘ��ԩ/7�~=�|lp;S�qbВ��s,�]��{�qOY	��/C&#g��/��B�O�:���4���:Iu�?3]��{�^��\0_����J���$��OxR@�]-=����C�Z3:.�Ʒyu8�ʋ�Z��U�!�gF(.����/�͟�����ꢜc�c�M����p�Aa����P�̜Z�N���-�0;ut[��N�^#��zˡF�Vd޹plT�٣�S�i�������ְԀ�
�Q��U;������C��)ۉ�_42{ķ>�.�qK'����R�!�3Qh�/1E0E�߀��z��7N����TT�͜+�m�Ֆc���D�=�k^ZXkj6���������<���2�����p��Jh?aʨ>0�^	�UǤ�$��\��Cz 4��b���~�v�&Zw�<�������&�}����ڶ@��|T��pZ���TS�C�����~Ð��_&l�0׉�p|ݎ�P£�>�uX���񻥚7��q��I����:� i�� ��2Z$☒h���.�(7?[b3��^3�+sNñ�K[��w�nVѩA��u��&���L�*���= F���)h�)FG���ڕ�5aMKl�E���B���������j'�Ik�α5qu+B�~D�3ˣ?�����V��:���˟���V��6��P�x47�j+��lܒ�ڑ�9������{���峴F���H���m�F��Ow��ވ���emM��C�3#�z*�]��'mō���C�@�7�grs|z��k\�0��ἤ��_9�,�5?��g	���5�O1[}���=�ް�Co�FJ�1�� �ǥ�ʪ�C	gVA��̣b��'�zO���֙�^�*Pp�����a�i�qҤ�ѻ�f6/��2#$#�1Q]x�UC�E�"MB$t�MUB�9C��	N#Sؗ�)a#~IT��C�����] �'E�bf9�Į�B;��[��h�	�,J�ЋP��V�ȐV7�����l�=�$���$���*s�gwN��
�$�[q�C;<~�t8��K��0xk>�s�O�c0���b}�sZ)���R����.�v����"]�q�:��ƫ�~/J�\S�����S٫'�j�A'x�8��u؞�>�b
�j ��ZՙY伆|e�:�P��~\�וb�4�������tn��LԳ�9�A�VM�B�<�5�</�eLᙵ���g�@����}9�*�23&���Z�|���;�2� +)(���+���%�{RX��/c<]�t'�d�E?*�ڴ��g�Ca;D �?L��
Y��>Ex��!�t>6�_��h<���J�~ �c?�#{H��ϧ%��`�c�/z�ZZ����q��qk|�\��Y�� 1$>��!d�������8YN��ݕ�/�c��]H��?��Vj�uø�}�mg�r��Tɻb�|�r�i���µ�ֹ=6m-k�
�ћx�m  ��UF�dO���Ip�ZD ���L�o�/�zW�a�nւ	�~@��+ph�@������6ށ���-��u��L�~���aD��0Ey2}���ߎ*�4ǈ�ٕ*^a��N�K�����#�&���de�j�� 9C��^}���^~Qb���! �o\a�ݯ��~r6�U1DC>�f�)%����$��ǘY/����v��s�7po��W��3���v��j93��`��aR��Vx��D��='�䎛XyD���'�!]� E�M����2W�tխ��5��^�{(��4Uph�Ѽz70=���E'�{�4���=��u�;0������� b�D[�Y�(��� �6��W���	�ј�/֡��������m�5-W��G����&XG'{�����S��:�����S���/Qhc��I���8
��k��p����E7FE�v2*�a����X&�O��ZnI�~��kM��0�[T��.���Y\��{���@*�;wCCW���X-WUI̺M���{�'_I6�2k��Go����}L+��;FxJ�|�K��cL�Q�FĐ��f�ֽ��Hb���L����,2#!
+�@#-��Z0!�*n:k���^�ߠj�K���-5FeQ������q�U��p{�V�Lo.l/	9���̯��1�a%��l�9:o����.ͻ��̽0��K��AML�-��2JVq�s��&�
�]?ZX^����V��2gmv��79�xQ����P���PV=��{I\�+n�D�)g٤�����G�9�A�O �k����Ǉ���/@���*��(�g�����Ǔ{b��=��moұߞ��X?r	��VWꣃ�xy�6�9�s���B����\��J��d�[����b(\�V�]g8G����9?���6Ti	�9�6w�_^v�|�^�(j	�ۤ�y+��O��ቱۚ�jV��	v�D�-���լ�b}N��C�hbyS�1����?Nz�t=��!��R�93�\�����[IݻS�|�g;��]WwE�'ibj��h���2��R�Oo���z�4N�vO�)߄�J��\~d+v;�p��}	�įwT�N��.@�T��#*��yC�
��Q@6�ٶ)�-I��*<nf��J���rV��$I�8J�0��>�
{6e^�&kw��ӛ�^�ǐ�q�J�T>�m��!$ү?%��m2}SĔ�9v�(r�܇+�B~P�k!'c` �T2d��*BR���e�˘�[n��/?���]��&�(�PV?<��:�����#����Z>>
�yiE�\3�������8-UAcE�.�G�hH���1�r<ǽ)D��:�#P'���^XR�_qxˢ�:����[��y��A�-F�-�-Q8��Fء/	*��mX�Lo�E���L���D^N>��M��U���-�8��i��=]��J�K3�/�{[�5�B�%vW$�=
���"�K�_��w����7W ���Զ��N(���E���L �I����f�������>Z��Q F��!��I+�q|�~�����' ;�<c%pNwը�1�>ቨ>v�H�(5��x3#���ĈP[�����PDo�\�v#Ƴv�D�y�/�8-;"������:�~̲��D~�}*����O�'ei�pY��@�4(���w�v+σ�u�*��s���� ��%ݝE��R6Z�CzV�?I�*r⬥!1d�-;�Z��xd��;4{�Q�N�v
�z O�W�1�V���N�?/R�)���U��G�u�N�Z��TL� �qcc�q�'��ʁ��ɉ�h�~��ʀ�=��"�|�T!�zp%k�&�ʇC�Ɂ1<��bd>��"D��C�SQ\�@H���,A�X����nV���Q,����Tq�@s �������b3�%?LR���h�&�B����i;��}K�邊yןE���t��;;m��a�^amH���Pr(,޷��C���I����o�0y������k�i#e�Υڍ'�DY��_�������X�,i~�ɩX�W�j3���d\�D�]����&s��J,	�y�A��qDԐh~	"G<���
�ݾ��a���k��z#���7ǮU����oP^4҅�g{���͙\���[/�ޗ��E����8ݪZ#�M
�0~2�96J0�^������n]�%lV�ѷ$3���?�L��1�d�3��*��:!��[�ǐ^i���+��`f�w�L�b��⁼��T�B�\�^nT��	�O(��7V��]��
f�/!��O4YS�9��]:�������^����&]�:�〡��,�z#�]@1E��9h�yv�)�`��m]�L7�k�O�<�/.^�#f�#Q����7�PH\����y�В��<,�(�_l�8�Eه�Y��ҁ@J�zaX�O�c�5щ�I��J�C
t�g�@#���K�Fy��0�Nn�Cm�>��y\���[;����ľ*����Ւ]�9���U���R�����b;x��·�oS� J�)f�\�D(#�B���Wo󶝹,��
K���u�!cϓ�� ��L��4��y_���� ;�0�-H�c#�ԃ�ˍ��~��D'I��t���Yu�'�.x �{�y��AW�C�L���V�3���	�^�ҙ^����I��a���� x)"4NqR�q{���!n�I*\ᥩB�=4�.bk{��t�O 8��ɥe�H�(A�� `��i��o��[�֒F����-%��;�����ā��B;D����p!]s�y���̀�G��9f��UFg�u�Y��37_�����.¿6ep=��x���Q����d�����x�SA.9���W!�n�L��.�	�I�}l�����CZ�UD��J��ZQ[1�Z4��8��pi9�|�#�=�(����"!ri>��9�S���v��ț)��ʓ#<���B�|�uj�0ݷ���%�>�@�:���d{=��`l.�CF�^y}�XTOؘc�6m<_��~��J��d	�l_2����Aytё'!��Un��E��쾥�%Nb�ȁ+֟�<R���)�+_gn���%�W��k����侼R�y��+�x�#+�������.��F,{���|軿�N�\X�Y���i�һ��Z!��p�1< ��/���0je�~������i���'�_���u�TT>Y�D�ꍉtv���Ԃ�/<aG��*�!�ք�DH��L�Oy��`d�
+�����Wɩh!o���(p�=7K�
�}�*���U������rT��tS� ,�sA����_�k�C��3ZI���Ҝ�J��]��z�;�.<�_>��AesdU�����2 ��H!�\��5�1�B�'o��z'nr����+��@#�m�[����fA��/�*�a8���dOE�K7��0,��z���^�i���w�f#��A]�Ja�\��
P�IȮ|A�[�pIl�au}��v {�Ay�"Cn�=�uT_�����
����JkK\+*I��B�[Ds�W9�~�C���$nA1�5�oG����=�
��vα��W�;�>�bZ�v���7yx��3E�oA?D�z~����vt�����L=?�	�<�(�ΐ�'�ڑ��!@3���q��}r��G��@��ĥ�0����V*��sUIB5aShe�piʔi�G�<��[/p�G��z#G]�G6���j����XON��ӏ��d��R4�Ro1��:u��q���5K��Re*f�W�]��Y�ʐ#d��ft�g����9҅�B����'1y�h7m�'Ac�����_�4�6�k|�k�O������ ���=
֕��E"��)��h`���å�-��G����0�-���a��T-0�������#�QL16�\((����# ��C��2`���� ��\�C/6Z6mި�E6;�]��o����ۛ,n�$���{Q#;�K�H�Kᡣ�j#�J��$�"�
��{Ȍ��̡�;n�H����Ř���e(�7��}��p(���X�)���jV�N����°X56�u�HB�Z1�Y��͇f̚�.�����mג���i�fc[��?�c�!�>F@��:j���s�@�)����̌6;V�7GG�J܉T�r�����%B7�Y@Gjԏϟ�%�|�|G�G;���1�g6$,��l�Gdd���DB*G2�5X�U�	rѲ7��J4�vy��M��#��3�|�RK/$Mf��S\q�LRPA��UkU����`�;��2"X��Ƭ�Y�-��g��Oi��8�\%�������q뻂�b��X�y��Fռ�PT�e.\:�v\+v<���]J'��C�I�^a�dO-���O���bt�<�$�ǀBg�t�I�����KC>Oh@�������P��爎눎瘎�J���X,���fWԲ�2gv�v���ѽQ�������3��`��
_eh/=�%���rՍ�ԗ�	s���:����Owع����(ȷ�e�T�t"�7�|�������dqx� ��xC��s:�hA��OiI����5&UV��አjo1ݮ��^	�m�S)�q���Y�*kk����A>�n�^\b��o�o �$�5���M�#��o�Z�i�J��**J� L��Uǯa�PH3�vSM��n(��I����F���]����$D�*:9�o�{O'���'�te:�<h�Z!Na�8�������(�q|�e��+?E2�0��;����8D�&ozm'Q���l�$�:$�X��>S 3؈4�{m=ۤ��a����c�b x�>"�C\��Sz��}����ꤑD3_�	�9�Ă@Br����`y��vI;*�A�w�/��6���w�NiYŀB��=��C�kQz��Qb�Y<?4�R�=@eql�՟�G#�W�f��`�-900+��T�%�D	�������I�=�LŜ)r�T0q3@g���DD���
�~����*Z����S%����Y�UF@�q++������p�fK��}�/�,Z�ւ�Ǉ
���<g��L��p�M_н�Q8���C �+ֳ�3�S�$r�@�%���Lਹ|���h
������i�a]�j	�JȐ%%�;���N2m��!���dXhhp��C��M��ޙH�#�w��l�{�k�cJ�3-�1�y�,�qa�zL�T/��b�G��ܢ|�M;gob`��SE�S�!_�m)\�1����l�m�lB>��u��h����\B�zAT�cZ�W����e�::��'cCC�����]J�{u%������'�01'�"k�����\!ބ
���׆jG�B"�9�C�@(&1%k~l���C|��*��� .�R���k}�PڔD�J�5�M�k��E�eY�����U;"�OD����1�6�Ep���Y�G�8��Q�ZB�`��A�m��̯x� �I1�1��9�����U���jD���7�ޙ0�S�Y��i�yL\;;��V�:!�Օ(h�aE'fs��*;��Cz(�Y�KBV���"*��:^�ڲ	Xጂ���z^R��Ĝгg�߉��3YW�F-����}!�u��B���I����e�||�y\A�B�.=ՉS�� ��-���zH_���8���wևNIGhꚚ�-b"���Q���f7Zl�=لYnY.�V���'[ �Ic�>���s>q��"��w�믨׈�'�6ۗMXdQ�%�f�9(>��}�ɘ+H��z\�O�$��x���6���~c�&!c�8H�0�1�I�ҕ�Uzp7�l�]8[���]�����60^;���]FQL�Q����d��A`�w�8�I!5�:
�^�[v�XV�[�#��!�4�T�ɲ�"۳2I�!�h
�X~X�7�?h���NǮ|���o y#��4�0��t߮*�6~��
{f�S�����$���������׼9�L&�A3U`�Ȑ�'�$�}�)٩��H(�tL�ژG���@,��'Թ+�*&5�Ӫ��ט�y;,d�.�Z+VB�0����NR}�&E�,	�O�6z���^[���ca*n�h~7gk�߰�O���/���cd�-�
���S-��V�_B��#U���ǀ�=�kO����|�WM�
���qV�n�5Ò|�ȼ_g��M��uֲS$����`���:���)+��3�P�Q�`��]�o�^uӈ��ӸJ��9G��|	�IH���jH#����ru�W��I^�H²�T��������\)r������^!KT�# �y��gtT�L�l(�����Pn���5Y s������vp���~
��ߍD� �e�6�j3 ��!H1��K:����B��o��Hi1�8�"x�fRЂ���j�l!}H��c����F��.��ԟCr<��!��9PQ?!��r��q�#"N��-������_G #���NU�dK�2��7����Z�:BTh�Qj����^�. &���ջ�<4:����<���uZ!�_'�^��^�k�/3�)*ۻ�E ���lb�ζ*"岗����f�檱܃x ���Ude ��t��ğ[~?�ڹt�:U�o��ؤE���9;\F����UQf
x��*L�?�^�w��6��.�Fa*�W-��T�V�.Qj����^���D{��j��ڸc}� 1Kj͠߸�D˃^�{U�0>��B�Ǌu��������=Y������ɶp�����;C�!�&Ls��^��L������6����^�2����4\^�l�`�ꎊeB
�_���I9�#�;+�c4����F�XH'����k�R`��g��;�zt���n���tF{ׅB@0�^�]�.��#�4������ƴ�� lM����b9%!&J ��\#�j�����do �i?��~P��/<{�.Qh$�CH&b@�����!ϼ}EYd�qK����}x#e\���d���!5 �q̫��V١(d#@9Ś1���)�fqU�	���_�r,�C�]R�T��Be\���o/��Y�Z�dk��F�4!e�o�ו��NB[��Ql�g�U��7���f�W�`)TkfI��(JW2�1����1��'䰢k�Ȣb�n ����%�g�����Z+��m)��&�;�E-��-��Z�I��mD�0KQ�.r%.R�v������C�-g�A�k|�@�r��8k\�ՠ�����I�au{i�]��]�]��z�M�@�?kF`����w b>6Z�(U��c����@ �d�R�H��a�.������:�s
ѥh�Ȱ"I"��p�4Ȯ�F���	(���摨u@B����wJR�p"`þ�@�T��PxBE�����|�=P��N�@wx����³Q�_�k�TI���_&�/~Y3M����_�ƯE@�U(�녉
m��D��D��m����,6�w% Lwt�_ɤr4Y����s/��nN*s<�N��2 ���P����"j�<�t�	��8��d����b��!6�7N�@��{�P�Mc#VHT��Nk[^�y!��2jw�P���o@�j�&9\���J����&���)�x�~g(�F�a�{����RwUHL/��Ф��������G��G��PI	�$låJs/^�'�I{���B3�����4����r�Qܳ!�V)�h)�B�-;�-�#>���l��R�@aZ�B�ut���T�x��p�#r7l��.͐PG\�G���Y�<C���~~�ϱDV�^�kזР�d�'/{N�hs�Iݧ��2���v��RMt�-2af��#�s���F	�S���25�-M@���\��7N3��>���䄯ͼ�b%t���3q7��/6pg�I-�徘!+�.��j2ey��G�U����%�G �5U��"
R(r'Q/9�?@�(IVI&D���3Z��iⓎ�zc�e�A!ޤ�W�o*������A�ʙ{\�T�?�[��o��I"���{4���odO��i�Q��.�<)�f�x����-y+$J6���Q�)��LN�I�QK��Y�D�=D�fkR�T~jv T��idL�1�TYr�vJ5��D q2�����t����I�R�Tj+�;oq3�҇CA�4L�#E�]��J�x8�y���l%��سR� y'}�H����)+�������+��:7W�$�">���H���N_��|s���W��Cb���Ϣ(�/)�=��]�@PvF�"�B;K��ӻny��D�����^FQ�2�Ϣk�����'ozזkR����Τz�{濫��h���<�}�8�[�L���3���m~l9�;)N���YbZ�d��8;���^��/�m��h�/�yu��J�k:h��&�x`�!��[�E�US<�.0�o��@@���tx�=�]kXC��i�m'�T#�z/9؉6��#	�*Q5g7%���|b�?"iE#�%�e��v�
B�d���m;��qv�rY�䛇�����DL)���C�[�E�}Q�Xt7HJ#%-()�tK��0��� ��H��-�Cw3t0�>��{�?���>��Zk�s�KX�$��HTg���y����0������9BJ�;�s��3X�w?�T8�d��\(��-a�D�LO�o!�O���/�C���M�1�8{/�L�;���&D����Ǫ��W:���UBBÍi
�)�H���dT@��Ǉk����[�=��ZX�Cm:�JS�(_�G���u���i�N��f������w˒��)���cX�v�a��YP���	��'��?oR��Z~�p�	o���4��i݈ꢞ���<�����] ���գ{��+�鞸qO�i��^,�c2{'|B�rL�����ǲ��d���
Y�G�����$�� �b�S
p���畉p�n�[�O˭�Xq�[_@c�J��f@��T��_�y\��Xe����v|g{�%��Q���Q���-+��e:sβ��R�ܷo��h�{��1��E�����t@4c�e֊ ���P�r_Y�Y��swm����U}ٲ\o��6O8�\E�E\��M�����T�e��u�}�ߠj���b�f�#��_�;8콄6�䜙�ˬ�>}����G�h�u��pzU�<��M�y���2v��P�&#����s��0Q�9a4#�D:�Kj���������W���N�>���!I�/�S�ѕx�]6jű)	�)~8����(s[��.�Qu����5 ��C��>�_�r�x�&�%U?�E"�4��#�X�pf[��h�~��i<�Q�8�X��L���a;�P�ebz��l^ͧ�>�����Q��~��B-5>7s�*�K����񰤻V)~���S�c�:ߧ�q=ky�5h�W)��d�½��4����������B� �r�sӹ@��r�i9	���H�����W��$ؙe^ę���E�Źs��-�3�2�	�6{��_��u����G�s�s��߅rH8��c;�5)r�+r�� +�i�����/0�y�9ʹ"����5���5�\.\���@�g�1�^l2ʣ�;{�Qf���>a�	2�@������hW�����H�Fnވ �|q*:�}/����͜��d�h�\h�;G(B��u�f�)��,����/k���`����	?��o�}�:����6�9܆ ����eM�=�|��O!���Y�M��~~qQ�[P�{��9��,|�k�V�x�v�AT��0H\�L>�`)��Aѫ��;	Uup�^څ��eoбa} x���9����B9ϓ�Z����
?�0A� 1�M�\U����7Ek��9lnm=uΞݮ4�t@���ɾ?R�`�%��r�s֏D��5(o�>��� |ڗ�Xq�>���yI�D ��O; Ҫ*K��Gg�� ����G�"7%b��`�1�-�'O���d
�u���{0ZNZwO3j�[=Uy�췥O�� ���e:)h�aST_<�	�k��+�bK6�:�3��X� ���7�(��!�Z�d���i
N��N�M��퍽�ّ�є����]�%G���=a��z�i�Љg�J�kQtBg�G��z�7�%b:[+<L��b�3uu��ޑ.�Ћ{@_�Ϊ���dw:�V5R�/�duq0�lC��&�!(�I��X
W��:<���&��F��$�W�#���p�T��)R<B�j�ծ�u�k-�n���[�S�Tě���f�6���������X��遨�_`�¥�ө����0��Ƕ�%C��,�V��=�j�۴�TCu{�����]�.��f������vZ�M�IvAԈ�^�A��=�J�;!���ug��w�cO5����殍��Ϟ���Jn�*N�)��쮢ff�_�S��*�W��.�Wʘ�Y��d�L!nS�ƪO�FKo,C��aLQl�a�Of�b�`��$��zZ+>tB~�l- >	a��ޗo6��0\�`cDz�]���B��]�F0&JRc�j�Ԣ��h1���z���U��#�w,��}�Y��d�o￐T�5<dy�X��-�&�hh$����h�y
��f3LU�����W�U~�ȔiDܮ�h�l�9��d4L�:�g=�z4똠����f�[y�0��1�T��Uh�*7o�]x�`�'D�ޘY*f����S=ܻ�T&�;������J��C 
yO):�Ϯco�`q��)�"1��$
^��uҡ�B�^��u���qyYĶ����BѼ-���&��;u��$�h�]T�s�d���b�Q���D�����3ۈW����	��uz���k
��z�lū��d�;���0p�/����,DہyB"��)���<G��fc㜡7�a�Ki���#s�O���(�� ��Х'�p{]�ȭ�y+Z��O�����^�l���Z���|'�p�[V&��0�鳶.*bleBx*�����'���x�_|�IG���ӑ	Vf���p�t�+��3�`�`O�.���@:�����ϫ�Y���&��gqz�C=L��5�#�m�b�K�&,�^y��f}� 񈘏� D���4)Hx�otS�|=��v7nӼ��5R$�p�{�t�F���@O�뼆�(Q�mbv�'�	Jl����	%�]2d��bƟ�|�	H3��^;(s+6�wطX������$զ��|e�>�n�XS������5���
��s�$�x���MCG]���nN 	���#�ڲ�#��$�����S���N�4Kp���tr�h8�Rh��2�)�^��wSk3(�Q�y���m�����-��Lr[4���m����ş��k��܁������Y � B���ݡ�N/�oJ�6Z.Ƞ��ƽ$f.�?��j<+�kT��6z�҈:KnKޠ��)
�6y�m����W���ʹ��=}�C2��Wר(Z��ՑN�M��dO�F,�`�L#�����G������/�����tK��E�	�vF:/ȏ9�����J*i;m��6�s����ڗ����)�=x�����E��f�PEٖ�����"���۫M$L�~�Y��{�g�~@9�@�������$d�#���;�Ki�̒:Q1J�x.K�ܩ��f�n���SO�&���TB�E��t���R�5%�H^�1�6Wd�U�j� )c,�s��|&N��<=�,�1���K����=�}�z�)?��Y�.9�%�M��f4 �E��j����x� =A�_�3&!/3V�+�I�y=ڢ�� �ɆJ�U�{.Wd57�5��3�����U�8���e6Y�#����gWBc���|=���������[�c����yAC\:�l��|���ny�.1��� ��u���� �^E=��ٹ��d%�1*:�}鿫���T��Z���b���kҥZ K�7�N�V��b����at���W��K�篧��˚��J�y��
���+�.�����"^V�ۧ�5r�K��F� ac�:��O9�M�F)l��l�7��~�³�����?m"���^P+�.�{N�qe��bF>�kI �V��/��?)�R�^>�@�7bgRA��8x(����B���Y���P����cYʊTp��Zn�%���+
&��t�1ōh4���!�h��a�j�Hŵd̐M�G�y����V1���!���7OZ�vv��ꛏ�D���Ku���W�;DV��uFM:��~�P� 8!)^tjF8����:6.C��g��0��&�R�T�Dw��#~�<B�_-�g^Q��]�3�RK�V��C���F���$����I�Zْ_�4��E�;��z������Tn�����@��>AK#�s��,i�����X��$�Epػ*�s��(�m�) �!ϣF.~?1�]Rh�_�U!�Ev;3���|�� Cݯb��_���o��)���흀Yi�;@�{��2�z�>y�Ө���׌�)K���f>Hb�3J� ��B�V5�����!�_Uþ�S(g��˒^�&��{����F�^�U���z�AC�1��Vm�<;M
��.6'����>�@Eބ�;{�z�$P�RnCͮ��+{6�O��WnR����5���tכr����}z�5qV�+X�2��ٷ
~5�$h��%���m�9H�Q�[����򣃁 "�uGЙΓЊe^�^-(���!��j䕋m�W#�}-������5z��"$�X߳Iګ~Z[�n
hW>7��-��_��߮��Ү��V���w9�0t�ӟ��Tt(����L��;�A�lH�KfV= ��[
��2��K��-�P��b��U��}ӷ�.�����D�\�y<�tq�Q􏃅hyц%��o�ރ�n73�6Yi��ʴ6��ܣ��R�So ��b��7��ĊTM#z�:f�	��ԝ��ˀB^&Վ];���y+$eTv=����yֹ^�7����[��KL"'Ϊ�������O��/RW
L�hﳬ�Z�j�D��h%JHm�娼��/�Vt��ndV:-��Xi.�i8���5a2��`���ƧY�)�����bq�v٪���TZ[�k'q9B	��͘�bY��B&l1U��Cc����PM	A�-����©�&�'�˪�۬PW�x]��8$�8È�e�*0�Z�����oo����;%�3�K	bk2c�o��r?�	�7x���T�S�	w���CP� ܁{���⵭G ��Q�Y�8}���ΰ����EGIź��bd̗l�u{����k����Kl�!)mR;
0�r�I%�>����N'�1�u���Ԝ2�+Q��s�<�ed��GY� ��a��8���#)��$WD��`ư����L����I=�j�.��3�B���(=?�B�+�ܹ�a}V��MrSn����ϫӆ�}�+C�_d[}$;Ӏ�:�r��`�#�(�[?E�o8����3K:�T�;$��}���g���Dg�Z��r���.�#<by�����0���8�C�OQ�u'��@���W;$���43�t��]�i�N�g����5��� �oz�d���^�eV��lL���Wo���HCO������~[In��Z�G��#�ETt>�
�;�k���ּ���(~X����|�\�H�w�E����8���-���v�ؓaVrFx�v�b'p�*�0��㗧ybYV��|�����H�J�i�L]�v��.��#�U����%�b�� ���E��.���R��(��x�)�{�����3�����m���EQ��z�P4�^̓r�\!,1վ�

�`�X���'����B��z���Yt�-�Et���Η���F�y�l��>���I/��r�Z�Ia�yf�H�^�u��d �|JE��1h6�
"G���?��l����z�I�	�u��z����t��<*�	�t�9��q^�O�Xe����W8�90��n~���zeA�0I|��eg���3��[�����Bi�&�W����cU\��	�#��9n�"�C��q�[d�7Y��K-�hB�-�:����y-T�V�s��Z�c��Gv���g�A�|���%vЉ��`B'���o?9�c!O�Zg�^SsNb�<�rTk�ٯj�ܴ%���ޤ��/k�
�P���M/��ק��+����G$��40����O�{ʼ:C˴����(���2��9��[�t'�{��\F�ot��H�$̝�Oo�긏
6�g��=u)����xJ���(iVS�
Q#��S��g�i�]��8�b�M���"���:���l��������ي��|׫�i�jTF�]2�O~ױ�����"h�o�	�v�n���R�"�?�8~�������>���~�ޗ뢗�AO%��y��\���R����nx6�vl�� �0IR��|"3|3�.՛�CR�\�o�Ʌ���v�Sx�V*�N����'C(�:�{0��#�%[�#s1:�ヂ�6�cL�h9Z��?8��ޘ���ֵ��-�?|�d�mpR�p�_)��5�37���ƥ��m^+�ܹ�s9��7�?�'^��ɂ�p�����D��>y5�)	.Iwk�kKn�K�KlsBI f]dG�9�-���HﲳԎ���]]�O9�*W{y4�:61~2�L�ī�3���ߤ������J	���c4�Y���&E��Y�*m xH)h,�;��?�K!���x.Zk�5�K��T���\&�J!Ixc,�,��;�l�C�&c��A�b$`���|��<����&9�nk6ۈ�&��g唙{L�LAa��5Ɠ�U�D� ���l�b���D��"�K����o�i�҅zN~��-3�חq�[�H�I�&�v!���6T�I��]d�O}	޳>�P�FD!�����A|��So߸��ȟ��Zŵ�\l9(�M�g�� ���d�7��)�i�[�0'm�pt?�*�� �`"��QZ��@	�Ʉߥ��(%D)F��W����oA�+�q�_7G�xd�;mVīNgԚ���e��:�܅��:�֪�o��S�;dN�}�G�|(���F�n�!�q���ef���is�񜵧��:����S��k�⼭S~�6p��h����W��i_��LUT��w�MS�Ȁ�������R�.��
�BF���]5ԫ��U?g�����K ���<�Z{�]d��}�V�kσ��T@��2�����?��B���>�|~��r���?��ә��s.9Ó/=/�/�
�a���Ήp�X��:�Յ�jll��.�<�ܳ�!�.�"l���-[s�j�n���:��s�������O�8��3Սႇ�k�6ǰt��X���&J�b,�[�W���SP������e���9���OÊz���t?d�U��T/Va]�s9�B\e�	��bI�UQ&�Wm3(� M�ۉ�������Έ�����*�z�2\hf=��2!*��}��_�x�ڠ�;:W��"��i�l��e?��KG������e2�Xg�6�ݮ?��}�p��E.��1����%���[��i� ظ)Z����V!�tc�e�<�7,*!�s19p!���q��α�p��p������|��K\iǳ��=��h!I�_���c"�
���h��H�z�޻��YR�����l�}�[�"��t���	�%Wq��3Rf�����X�zq�9�5��	����/Ua"�}ڵ3_ׄg��:39'��_n�F߾�NS�)����ij�gU�{Dr����M�l~9��?�����&Z�|S������*���W���}����YEH���<}���~# w�	A�%);Fm٩Ȳ�i�����{��3�+���ܭf�&����-�X���{���+B���~��f�PlWC �#i�O�`���?���p��e����j�+��M!�n�6+��2˖����9������\K�)d�e|�!FH!���u��"�ip�e���x@���g��ڧ�I�q!y7e�ޥQ�WE�+C�-��v�6��T�8��zb�hMD�Նy��|�(� ���0i$<I0/�r��$J���8��ٌ>�R�[M2�i��y����~H�\�F�PQ����������>�$�X�,tM0�	��n��G��0��[�HI����r��J��"�̿H;ȡ���ķe¤�*M/�_03��%J�>�o""��vȜW�V���AP���� ə�űߩ$x�B�6 ����WД.nۡ&0')K�ӕ�
�$Z��K�t����J?�A���w��&G������<� ���Y
� �ÿj��@� �����;��G�pďqc:�̉ƅ�l��V��iv+������Ռ��������
\�Sau�3�.�!~d������S�B�]'�G���,��4�sH�ď�`�s�ml��SP!�i��'yynU���]`�[��������)��D���r���W��yl3!K��!��Fq�r����b���ݝ�T�m<��>�GuҨ�g}��V�'�H��q٤}�3]�\�ĲyEݛז�!I�s�	O؍q�%�h���Zr�V�=/�Ns��1�.l;=�2��d����㌷m��L[�?��ꑬn�Kw�IP	�RBü�md9����x{��&�w�-��)�؆V&�"�#{�j�%ܤ��l>��$�tz<Sm��H �x�~\"�Ka{�����5���ܯ��%My9��ʹ�=�����m鑋�4[��WG����������<�3�d�Gnk[)R(���k�s���[�~͒��8���-�a�
 %��j �5?:���$!l"�z�myv�˞�>y�']�xT�v��lţ6��L31%�bC*F��Y�=M�.VS���xN�*���%�%��}B��2� ���M�7[mW��T�B� CQ�㖅�&�hrW��D�.z~U�{�e���tF3u��'��xaTM3%���+����Sr�b­�^"���y�k�`%�z]�H�a�]���Wm��8&H�Wg�O$XxM�7��p\(i��v�ےfS�s��|\qHN����gc���v���Y�9����<��1k�x/1��d��a�un���3��y>�_�j��"��h�0Gl���8�U���.w�y��NA�Ŗ� �����h?k��z=��̘H��������Mr�4�v �޻�v��{��T��G6[���������8nv�=�
�c�V$}��P��������ӛ�R���W�Ѧ_"�lD���a_�ۥ9�M��c��)2M��q�VH��� `3�� ���*c�&�' de��+3�-��Ρq��� I�1.6�M�r�gd�N�4�>���5{��8'8�t�۟n��%ya�O9��eT��I�42�P�\ke���~������8�nC�Q{-~"R� )�C`��(��2,	圯��y��*����\��F�J2���r��}�'�]q�l�ֵ~�����K�X��t��e�'D.p 0�#��du�8Imn���	(r��'J��I���g,H2W@E/5��qȂP.��>"�о���*{�pJ��4^C��K�0u=����IHa@������\俰�x8��;i6�|%x�5V̭���h��F.��[o��M��%�mc	5[�8���6hH	���2�$��X7f�Tr5 ��i�F��9�C`���n�����vb�c���y�re5���~���7:=�s�FH��p3ǔ=־��"Hm� �ԃ<��=��lX�Y�pL����o�`�C�=or�M�blU{=Iu�<ֻd"(��>i��]���H����.1,Dї��9�B�Ӏ=nQ��A/�ظ���f���R_�a}���T_��{B����1�G���R|K\�d�f���	���t(c#�� b��*G��]}�'U�~>Kҩ%���w�r�s8��q
a�i����CҮuQ�*/�����k|m��+���^O/k����xy�x�w��`��=Z�)�����Χ�-w����_��k�8��'d���ujiW��}���C���������í*�K�+DQ�������3���R5�<�rF���V��_�f����倲Y�������D�o�<�̳`��GrC��+���2+U�Ƿ�[?��x��m>�e�+�|�P��c{F�3��f"���8���tji��&�޻F����}B~�+_X��T��f�i�/�4��?�D,d��>���n:7i
ӫ���m��ִK���q��3���Z�.2�hu��y����`(c��W���ݶ�ߜ����|��>��5�ඁ _*B'= 5s��I-is�nF�Bn��	I���1GG��Wl�ƁI�7�E��0c�{wf��u�u��	�C+<�{��v�����k����9e���-&s���~(�FʹI����$�_K��@���=�5����Ls/���Z�)쫦�U�}a�
^��-��2�Lٳ��@����wz�ę�[�~�h�.hA�Vt��4�7�P�������Ϋ5!�3�����q�@44��)�� ��<�oC��i�I/w���Q���c[L�	����M{W��^i�9�rLW�Y�|�T�ۄ|�� |��us�+J/bh%�QN��Ba�/�aD��Q.81M�S��Y��"V���/�X�M/�����
����KF�hy������ ���hN��W�\�H���`��1�Na�����������n�@6�8��5�7؁~XF(�i��d��{̏I�M�����Te����{���jG-��+ �F#{�5��Ch��w��OE����o]��/���L.5AdX�9�����g�Sg��Nٞ�nce���F�A��4��t����Wyw���N�;����x0�u#�:�N�ڲ%���Ѯ��97�h�)�Pr
�K8�TUТ�+RCsV�/��LW��Ɠ�4�X�\��ڻu�l%]�5�®ʹ��~n���ƼΦ�R:�h�DiR�gÚ��_ƕm�t�^胊�Rs���:�H��g��L�+,���c%t.k�)c;�	� �͒�[��������+A�E�9���h���`pV�D�4}�Յ2�ALX\* >̌IB�M�3��p�Ŧ]T���5q5
�vӊ�T���Fv>����v�B,��M�ҙ�K���鶽ܘ|8�4�hG�M.�u�k2G�b�v�c�:�]���hȯv��9��G���P�^ԍ�cE~&ʓ�mS4�OT��6�2��Av���������)����!(O2-\�Nb:k��y��H�����y*x�yG4|oy��7�sݟt�����TƐ�z�B�y���$(���t���OR����]��GH��~f���;�`ΕVM���!�|H�\�Wn��Z�'�^Һ%�X>�.p�����Z�zm��eN���#q����.��~l��Ua]�P�r���	|��SZ;rW֗I;��}d���!a��R�kh-�՛�1/	�B��]�7%�ll��b��dI�@V��@vKESO+��Tm�}�k)�Ȱ���qͣ�q茌�VS�B<�\���R/���qD��ˉ�Ӻ�ڽ��E;��z����Q3���	 ��`�-��/��T"YZ��G![���L4�z��ѿ��a�7�-5�X��%: �t��l"H|��p�_Tp�t�'w.��l�Ye���C0�3:������E��;�Y��z����_�XN���u>��5v��C��_�k�:by��g����+��L[>�zn,l����$z���t�N�+}�0L�0�+���F�t����u�!\���tm�B)n�Jebe�߄�.�|*x�N��n���z"rHUbNT�i�;U5�����xG�-�w����m���I�����7��e����O�9�M�	�F�<6�ŗ\�Ҧ�)�!Iب�Ô���C�|�]�
�;��E���;��D+��95d������n���318�ihO��͒�pR:?�5-�k��6*禝$�Vnв�$��_tn�����q�*��p���r$Y��R�"��ˊ�U3����5�Q
_��X���9�+���	p\�p��$~��E	Wnyԛ��l�yS$~�~"/�aȰ��?��Dʶ�8]���FB��=6V ��� ���k��;����g��3i�4�0Q�>^?R�s��l����p��bf�vپ�p���u$	���:v�q�W����5)p�|����m;�2����>�_�4ꍦ�n8�]��S_���v��Q�U6G1R*y��c޸�	p>j�Q摒T\��8PGE�a��xϬ/R�c��	C��U4K1*bs�ǡH	��.��Ѻ�G�Ϥ/Hq�]��"��X�]����I��Ӓ���0�7�b6~��SBI7Q&>s��ӕxs$L�_��������c���,��Z�7$��ڥ��twM"#�b��;�q0D֡�dd������s��4�'��R�2/i�co����o����G�!�^��^Tjl15��`�����u��b�	ɯ������g��	+���1��>���/3�w_
��E��2%P���_�q���pw��������up���,�g��� ���CJ�.�:�j�<��ʀ�k�m�ӁԎ�)�k�q���h��m���%�:_,��p��'y��?N�t��)Mpm�e�[̇�_��>@�*76�b��&��l�I�m���5���u�8?i�����	/�%1���9Tz��`0��|
�Hk�2g6�떦��c�x������������ϞM̏dCx2v.[2�ZL3׶Cp.��Fht����^aY�>�A����w� �s���V��͙��s��R�asc
'�nL5�N�c��8��ςL����#��FS�^}����P��U�;=�;9=����2��B/��/�0b$�԰˒n��q�|$~/�N��qY9�%io1``ȍVR��X��y�Ȥ<�䖇�I��ŵ�n�
�c�i�:T3y��į�r�,Z�,�����LJ[��R;��l����M�E�ɡ��-ٮ�~�},���i�g�4�?f���|p?�whW�k�'��wŲ���><v�s�u�+������������CfЦp��{np��#��IaR�O+&����%�D��6ϖ�
��w[գ�+���N"{�lP�ӱS�g�Y�D�|���P2yӔ�]#�n��+s3�b���+��*��
�X��m?�O[�<�o�6��j:�!�&��k��z!��Q'�D�_�2�>))+Af��B]t>+kd����"J�3��3��$�z�A�+�lc��o}�X���e���ZV�x� iOqhT-A�$�ֿ�s3�����9#Zh�>���x/�8���p��3n�"tB�Fn�p� h��ئ�6ȼe�M�3E�r���/�w�k���y�/ Q�sڟؖG�9���/���4����&��Y�j6�fa\�؏N+��߿��JOv@��B�q~���y���쁉� ƀ㦒���ꐒ��N�f��>T�ȀmhV�s,�<�� �6�Mew��%��Y�����Ʒx�|��k���7�ژ����R����g]�q�����|~�P�]����$�^�E��{k��o*���A�R��ɗ�W�R����#��Do7��<�8"�$��8���}���\��>��L��rlߑ���s2<N�n��kV��(�j�
d�x;)bR�%1�>������&���!T)�f<�P�j�7tq�xK�ejp�i��2N�l{:�	����R����vH�a���i�Rqpk_���X`�-nfi�c�a,�	��<��.�쳽��=oK#�?_��4�T�����@o���zS8�qǭ�f����4%�KϺ��O,���a�� n�Fu���"鉊�:X��V��_L>p4m�˜é�L_i��!�"�[��ɛ}i���r5�IC�NM��{)MS�����e].F�r���hh6��$�f����f��z�3uE��j�YQ~J���+�*w$�������������uvq��0���<��Od;N�-x��x�/��	��;�ܙq=�6Dy�����mv �����(��T{jO�4�/W��]���K;��Un�l}#���	��S����-����V��MdC����;�Y��o�
�Uun�(��:����c�?3���s�5�[ʋ\Ba�'���i(�C޷5�̂i���?W��L�OBᗙ��t��,�ݟ@K>�޿���)����^c��%�VvoVG���,��]b�����x ���|���8�kC����Q"�I���=oɰh��{�dj�֮�(�r�h3�&����vb���U�㛎S��#��7@�ѩi"�5"������9Ξ>���(�5mo-��<���6#*u��2ތS��z�%]��q�}�	���~5����+^<h=}����|�O2SP3*�!S��d��r�RR=k�V�c�Q��hk`��f���fq@��et���p��F�6�V�n����X��K�v��0��e���e�A��Gq#WB�Io1�cv}��:�k�6��n�Ȼ-��E��\��PEŕH]�oL��3���G)��m�V�uW���Co�k���b� ���TW��ɿ���ıK�.p�4n}'��@��������T��wu�8�7��f|F�qn�r\z{:I�h<l�����|��]����@N-�I�f�>�mbu�kq"�Z�A�"U|���I[��&
6f�����?2`��PB�D�tx_�YS�`�%����D�G�|���3��2��򋕹�xW�(N����m��\2�=.��>����3���Lq�s�)m
�j��X�՝˚��Z��hA#�x3�\��I)�19��3��.�J�af���3��	ق�aMF��4��a��T��-�aY'r�c$�s�£߸Atߞ7~��'_����W_$&l<��v����c��f�ӊ�t</��KRF��m��O��<䕊B%�2$Pj��o:uڧD������,�1�S�+�{}�	��
��R���r<`�J����~� z{������*�969�iU������Y�d�}�?��I4�� �U,H�k�i�ژv_T�^��2FjI�����>�@�]3j]�}�z���"�Wq�V>�4��E>f�m�
�czV�"쀳�'�u[�}ékgG=�O�Z�³��&g?>��:�yJl4�m�pP�6u�B�ym�My0��}�0�ۍ�'�a�ϓ�W�mpIɣ=��R�b��fmt3}���w܈�Y�2�	;fYP�KYü�!�OY�I�b.�����g��jY��l���ni<q]��ƛ�����Zؗ�u�z*���`��c'(`�ʷ�o�#�aY�	�V�I���������%&��E��g�f�"�w�p'����5[�	�/�;�R�I�3��2f�7@)��j�>;3
�xލ4�����<_��#��XA��kS�C�d���R�e�Xl�H~&��-����QA��e׻QP�>0�xϡߺ�x]�a�.��P|��H_R�ae�z��pe�S��6K���x��la8���6�&��X���%WL*T���%_�+����}��ղ,��A�!f"ʾ
E�����T86��>���N�*�0�:kh�D�]�(D
��i�Ƚ_�n?}��r�/� ]�W�f=p��鉇��{�\��
G�/b��}wgE��+1JӘ����|�2J�L3n��#������a��j��sY�
pd��������0𮂾ˌ8�e5=�j��7�>�,D� gї{���N����ў�A�z>`�rdt����(�@���ƞ�D�K�ޥҶ��G���<���$s����5.���v�ݝ�R>9Ȫ���g��g��c���)�6$�E���|�h��z���!$����<z���l����4�ı��#|�����S�m���Q�/�4�_�ʜ���l��\Ĉ�k�}j<iik���R�1<#��ux]o��=�͆Ȼ�B�:%9h���������-��By�oR��U�-����<�ł��P�-�ȗ��j��0�����ȍrׇ�ذ9-�K�}M���R���'Q�3����/��򂣓��8Mz��]7QF�s�V�]�>S��z� �'���^��4 ?I��/��?U�,/��L���n�`�����|�REy-_��9^��Fuݓ��E�*A��k�V6ԕ�Zib�b0���ҭ�4|�����+��u��W4ft�L1�]Gv�}�]p�[�R	��� ��v��6˨=���ZH��>5�&��������B�v�d�Ƀ1|���elmB!��\$t�eM���������^�G�Ԑ���
��:�.�zG*�Z��dm��e����^��p��e���F���c�s�קM�=��|���>;" ��?�15P� x�./>$�����8��
�6���s*X��)��u[�zGc����B?U��C�?7d,O�k�{��N��;R�]{7EՈ�2Ծ��b��P�y����ȧ��ɏ��g1�ы�e�j+|o�i�2�#�I�r_6�#�Wh����*>OuF�%#��k09����P.��`)ީ� ��3���f�(���*ڮ���!���+�&	y|���3yD�!p1��݉��M�P)���U�3jwP^���K��-�0@d�UvY�q� �!�&F�h�\��e��	A}�&D���?d��#�f�}J�㖬��Q��A��Z2B�Xd���=��X�I���Qrw�]�+��<`s6�?�l#��:r�O\�o���_����T��F��sg���w;k9��!���)�~J"�Đ�CU7{�A@���nv�&ew�L�+R�7��Ih����F$�� ���w�y���@ Lj�dk61Q����a��B�}�L�|ki�.1��M1
��+x ҅n� �H1���@�n6��F;����b���<��m���s�hBL������
�o�$ �y�2G���������y
Q!#,�n)�U
t�_�k'd��}��pF��O��I�3��t�?��>� Z�H�7����)�/]�}B�&���H�?��
�@x�P�;t�i�u=��ox�՝*����?br����&&�{vOJ�UF�x.�v��Y�c����
�G�##��! :�Ț�Dп%y�G|�=��{4����s�Z�AN���N#
i �����%c���O��]�S,�"�X���5�Z.�y��ڥ_J"��U$拏U;���L���= "���J4�GE�M���<�S//˅�~tm��TM��ٍ�/^x��*}�5�Cs�r��)���o�8��U:�p[\	�S�H-��vˋ��c�#�S��>��|�������6�
��y�A�>�P)��<����k�b Տ1o�b�㤯���w���[,�vC�r#!����g"�f�O�@�~O��T�PU��Jww���� R""-��;DZ:�I�N��.���\J�޹����7o�aƙ}ώ�Yk}>kﳏ�ėOh����|~d�����f��n�5V��H|U���:^}������T�N� AU�c�2u���ڃ���;��r�q�ym��Ҡ�2�XSp>�9�S�z<��Ip��7|�y����I$ؑ�����T��K@���*���'���@i.Ћ��7�!���7̑}�H���2���3S>'*H�����{7�Q���:o��?���]�v?��qG�`; ��R|�=��Rՙ�����(���Q�3�쒃CB§j�'�^r�`����D+S���_A��iǳr��������~�{��D}:l�;�$�U4?T��9���g��8���GS� ��_��HU���r��0Z���_���� �fj��2[$��{� ��3��T����q�D�즐*[dIˀ����)%��ˣ?Ƅ^Χ�j6�A! ��x���h���҈Pv���Խz;�a�1A����aHx�:B�U}|��^95	��f���D�K�	0S�+��!l�m��N�3t�5�����%�&�^�=�TϖJ���ֻ�仙��<�i6��ϝ�k��Ó�ێ������9w�o��}'-m�5�j�&UƁ@��w�R��e4 	�D��Z݆<u���FO�zVUc#��`0py���F�X������d�Y��­�c�؎��ˊR� x6�-��' X@���v��7C��Re�_��z����;�;����s'�������/7�ޱ9��lC@�]�RlkG}�{�0BO�{�,����cS��^Q�n��*1d�\�@�t�:k|��%Qb>M���T;��]]�U�8Ó��F�����	@�R8���o?�!��c�K�K��7b�ϻ�|h
���-t�j��5�]|2��әv���q�W�z���);�3���"��ɺ�^Y"��oR=�X���4�*�๛����B��S|}��DjE�	jc<��x>S���x��&g���ȢFX�<��V�c�_�)�ٟeEg{�_��2���ª��v΢m���������]eT�ѡR��ҙ��b���~�����~���P���x�F���7���/	���'��2���'��4h����{����&�lx���	xj��$,^�Q+rH��䕼[G��Ʒ�mj�@�dq�*���j5����2��'���}�nw� D];�L�|f�'�����C{��_9�ѯ�0B]s=�Sqy"l��e��ne��CՇ╍�2�� D�
u	^���^�wa~��x�K7����ʔz5��ڮ����-�v��DۑJ������U�tzl�Z��#jp̃<�q5n76`Y"#X��&��0��4�,#:�];�uSG��o�������Tq�Dd�rB_�	k�2��? ��(Zm����Zq��8V����3�9�i�gcuR���Zc��X��!gs�Z�]D�7}-F@�Kl����,�u�d��$�ըV&��,���N�.��#�I�{����f``��b��ݕ%*Y����p��[���@A/%��{z��齓�$i�lG3�e*��u+Cm�5�Z�P8��ǭ���{CÆ�]�֝K�������Ʊ�蓗63&�p�r��53����<�9�F�,#*̓�-3/�b��9�lk6i��|/��Z�":��ya�Xe
�j"Rr\�95"|�����94��M�(�Ff�u�\�鋞�SxB���y��+��_��R[]O�|�KG�BVե�E�&���>�l)��ky��@�ы�(� )3���H��U95�Od�=�`:s�R���m�
�ra?:�X�E~�~��P#��K~��iw������'Kچ��Y��=�S���U�����>�� }�m%�2j��rNo�eH�����F�*��`���:�	

� O���Z:�b?�ɒ�^A����x�h��K�;:���~!���^�GM�}��J��a�2���ճ?�\�J��N�k�a�~��1�R G�ݎ�&�j[[�R�F �묅�KeX�J/9�vV���жX��/Pqw�iA@�ju9Ȍz/���o��'�NX)��p���!�.}�艹�BiT�uT�Z����Ͳ�	,��A�gm�z��>"zU�Jbve^n/L�<�qp"��l��s-v<��kR�p��i#��j�H(��E�Y8z(A:�8�����Y  ���� A�Z����n+���3� �S�]�qy��]�qΈt��B#ʿ��<�rct��F������v]�&��XZ�ř�ńҜ]5j�F]=��"�$�����L�ղܱw8s)uu��h��eCl{��b�\�!�L����_�r��\�����b��Ƽ����]b��>hke�~�?0]�<ZE��-�?��ogT$�b��aa�n/��K��@���{�C���������vZ�ŴuB:�|�\BHw>v�UR�c8h����Ng��fcپ����N�T>A�b_H|Vqm�@ާ��و��}ҋ��jܠB�k�s�"��c��+.HD�q�9�6r~ ��p��I�16����o�1�X
� �6�ٝ�g	��d� �}|�����4������xM ���~Ů1`3HapT(�S1j���k}^ݦ��VW��DJ�=io
7onh��'2��-l[�t�1֛��5<�ڈ�*� �$:ڝ ��ޫ�]ڊ�ր��3J�̴^�Ӿ�4�����^�����gw�J�`���J�KG�J��V3���@��+����u�f��d�E�mlN�G/�9aH���>y2C澂?b��K�xe� $�[L�+O�э��~Dc4D�WG�0odx��.J�0�	�O� �[% ?P��߀��P�a\�_���*S����w��o]c 8�c-�M����0���'e��1tz����J��㩖�|�H.�V�7癩`���e�-��/�H#&L]����|pO�3���|����8��Ԉv	�㟌�}��F5��/Qs�=5ט� ���� M�a2%�˃S��8����n�E���̽�w�!�*��'$f;#���c�Ly�=��YQ9͸��5�}
�|2G���$���=�=���k^�p�wZ��_���hX����b���;����b�x��Y���3��@��'�j�~���0�(i ��;�Ѷ[Yd�d����c�ei3������PyB�"|[~��Id^ �F>}(|��~F�6)�M�k ��c��3�h}�w�cs�p����k�R\�:U�b�/�O!#�W;�F�5�fZ�m�U�ʮ %��;�.��?1Cb���� V�Đ�v�]��.�˱	x[��pc�Y+x>f��M�అ $ ���`)���W5����a�$.��M�^��H��4���7vx�Tr`ч�y��j!|�v:k�v�R'��^��NED�1d(�����w�}��]��C&���,���`�5�[#?�Ɂ�3�0BQ��zx�����a#/��,�1� �d�w�g�P!��pK����A[�ʳ-������G2�L@GdTN�$Ⱆ��0a�m~/�#�0����,m	ދ�D�l�s�n�$[D\�>̋��o��w�t���e���5�ց���?t}L�%D��9�v�L@8۟$s�;aD�tԹ^�ę�Փ�M�p.�>�T�d��\f�&pTV��F��+�lR���M:�8�S��} f*��#ry��ϓ�yL�N%Ӈ����x�H��# ?�6�
�}ؓٛ8����`FI(�-Wޮ�}4�7䏃@�1�h�W��5�r�F� :�#���2��I�2����t�ƍB���eg�����m���^�v�����k����#�o��͗��g�mU���'��)�]�
�K���7%��I��5���a8�,90@��΄�Iʽ��\��fߩ����Z������~���M�MJ"q�	}��0i�W����8�1$���
0�4��rE��0l$w��3ev���۲�����v����0�芾�S�ޘ��9Ğm�F��PYEd.S��8�`�%����z)m��Ƃ�/��x~:M4�)ݕu��a�����p�z)+@�&���V�]�ۯo�9���3:�-+�	s6{�l�O��Xz�$�#��Pv�vU�G�KY��}����;/N�mi� �y['���{|��D5$�{.�
K�k)�1]��,����-!T$���0�X3P("������h}�5*V�J�i���{+:��/FSPdJi{;)C'|�y����F��Q���ꄍȢ��$HF���y�|�A���Qc��B�hM>�Q�"ڵ
�����P�����	�
s. �4t�!�����,����~��3�?���
�'u&��{��9�����7��qMed����1��S���Wl�k;� �R����<��D^^���* ̔����-/�).�X�����f5�.V��wi����Xچ�/��x�b�yŠ|]����pq.PQ�5��i ��1�L�ͅ�>g�n�Ã��uf4� =�F_��{Z��6��$�u��*�;v{��}��Ӽ��7��z���bԺ>~�2J��x��m���%x�����2Vl-����yA��c�7փ޹KQ	�A��D>��9�S��T)4�DJx�2#6UKn)��	6
���z�WБ'��v�l�?pI�Գ���*�;���減=KTJ�?�����gӔ*��R���6�y��6�U��C�u�����jG��P5si��i;�1���.
����)F��zx����bZ�Tnq@0�aw�\��2��!e�!�v�SL
��."8>^ӷ��=e²քgO��vc$���!���'���##u���Cy����+(�_<��=�e��@Ν�x�BTG�T\�̣�b�g^�䜁����L!�&���p�Uj�#ut�3GL�kNŌy �G��^�GC���:��,IF�X�g����[���c^8<�/%�M)�Qq^��w�`؈����\��SV�r�;nøߛ_p(W�yF���Y��m����S���(̍b�ďQ��vk���� -��݋�w������qF޷�,RCk~Շ����El:�|�\5Lt��cc)|�mh��T(��,��$�ܵ�ˇ;g��� �M�{Peѕ� Hdj��+@x�p
(�$�nQq��!ŎQO�UFLǿ�V�彖}+��bwIde.�'t!�p�l�ܹ�=RSs߆�C�~��{Lr���f!V��87)��64�UWd	C�~T~eҊ��'#���^=������=�!���/�g���U��F#�X!b�������h���K,��de�}�ȯ�.n���D>�Z�9�a;�ZSĆ�A0 �V/��R{��x�R��[��y�.#G#1Ֆ&��e��UU�})����֥*�4���٦�F�d[^��s��
�ҋ�傇&�?pT��(T;:�K���Ө���H�E XF�v4@6����㗗��F���s#q���d��P����=J�by/͌p��]B�¦�����t��1��^�7 ['�^4a@���/��,�Ml��/T��ܯ��-�"���n�&Z��&%��%^v�F��(��b�g�V�d�w�zO�W\r8��������S��}1ެ�A��F0����>[�G��dZ]����Z4伣U���f$���ejn���	uNcQ���ώ]k���E�xJ����*��\
A�/�5�@n��fbُO�{����Ǿ3Ŝ:���1����M.�,���� ��o��k{�n
��sT8�]�ۧ�]�}[߬�F+���hU�`\|-����`ťSo|��T����`n�3E�l�+��\F�����T��˵��>=�Vibm͸X؋H�+5	���| n��A�V��~�ؓμ�x�`.�5@���� �4�*����9tHJ#O�`��7����̚bқ�J}��'�mvb�Tk\�B_����T(1��͚��o�~�,L_: "���}~Z�9ѣ��V��d�����G�� �wBM_W��8�!���.ms��&7���?T+�?��}]�,FǙ4�D�;��ͫs&��_=���By-��m\��c�x`ol��8C��I�s�u�X�C�o�^D�^�5�P0�����z��)C*�eJ�P�͊Z���N�S��DC7�����f烺�U�V�{L�h"dp�����(������YV;xŎ}�I��y�:k�<F���8bް��0�0]9R�+�-��<����8Q{��O'I��hۯ,��	�!�E��^^�nJ�T]V�ϛ���_������=�|��6����jVbV��%��BJOr��D�	��K��>�E�?�{�.(x����ח� �i��ڐt�|
��e�GE�d�sy�\��;� ��)Nq�?��N�����ܞ7�����0J�?<^g3�l1�ҝ]�x��48OV���^+���<��wtT�N�� ����qF	��� ?�%_��˂BG9��:\i�~(�~�ݳZiq�ʧ>�NHZ���hqGE�R�N0GiQ#}Ztc��H��Ώ\A���sԁUF�|�(]GE�/n�ߙ��4����0i�����ƧXgK�d���d��w�bU�)���]y����B�q�ʢ衭�_�q�'���`l@c��b31l\ӕ>+���G펉�O�&�6zx��r�����:ݒNj��w���8ۻ���]�����f��ӔF�OR՛;oE`(�J#To�����|,խ��#�d_�~<|���/K����Ե��1��ݔ�n���6}�ߪ�)�C�oC��te�$�V�&�]P��7}���¼9�!����Z*\ p��y,��
�uWam�6��4iPG�lZ���pسu9��ލw�Tqm�d��g(��U�q����^N�:���q���o�����j�@=^����d�������ݢ��ߌ� f��ߎA�d;���Y>���ڐ9���V2��@�@N�tD��d|.����HJ�CG�������[��[t��݄ Ճ ㅓE/�c�yZV8|��9#i�?��Ҍm_����k���J��( P����.��W�~����Ɇ��<;��nd6�P��6�V6�T�~~�D���'c`��}��{�M�
Z�t�,��o����_�*xiu�ұ�B��{-q}�E�ߦ����D+a@�HJ�]�����޼CO�mYt�4~C���7���A%�y��5	ߪ�Щm,�`���۟񷟌\���󥮙�������Kg�}��6�,���O�R�3ʮS�K�Z�N��1
xG<7����a��4c1Cm�@�rm���yG县�Z��j��K���/��%�˳�`A`���v���<Ðfo@�����̿Ώ��TF����8�*n9G�c#�1OP?��F)��&s+O+I5.���
[������t�JfU��n};��m�$��������V2�j*�{��Uk@rw6C���1 "�rKI�,�l��u����a&���m�	���O_n�2����?Ո<���ӗX��[x�6l�M�C�|��K�V�-�;�V�}s��W�䐅�,4 g�������kq�k�8�c��8l�L_��5��$�K�Z���ɿ����bU��[���.����ꘐk�d=�eM|��s1Dd��+����>���O/�%�c��)�o�� �t����s=�:�����-D���׳9��]Y�P�c?��9`S����)�*���)���-��ݨ�+����rӇ��¼�PG�#�c����w�^����ڥ����{�l�ը)~Ȋ��(b�	 ��/K��9���0���ɭ=?�����s��Շ�1��?��)6¨ٙ6�/3-�d��w��y��^ 'Ӱ��x�������� ���nE���ƀ�U��a����P�|�?PK~��R){;��0ds�����B ��P%�4_�N��.}�Z��gg� �a+�5�	v�u+^z]�A�W�@p�9��-�i�oƺ��H~y�z3=R&P�[�kW�T�(U�q�6-[���]xy��1!. �R�����'��j��> �;y'%ޡ��L���
�#���v�����^�x>�[NW�x�d$h��� �����_ڛ��mժ
Ŵ�E�Z�9������j�Ƕ�^�ӛx�\�)Mn@h*3��b""-~ﳚ9�F�'����״��|�W�j�*�#{�o?}o�� �~Zl�e��"����`1�Jq�	!�
 �J,�#6���P�lBب�[���w��|�-�J/5�Ũ� k#ޚ�g�Sm�jz_���S����t�F���ȯ���1�|��}�}3�.�T���P|�DN�-�9���ˈ�g9��F+�n��p��^�����S�ÁP ��jk��#F~ ��S�鴗�m-�WQ�	���τ�G�isg-Y�+2���R�~'����i��-��q\4�&h'cyc{��N�~�V��4��ۏ�[�e�"Wü�{BQQ�v�Јx��Q|��G�!�Z+�EE�'|�� �넙��ϘSF��t��ÿ�g���k���02�Lavj6�ޛ%:ig����)������^w�dę� ��L��;ho����+	�yPh>GS�[�b@�i�%���������AT/>�}��2�/���#���*�f�ax�FR�l�y�����}i>R|��>t���t�̳:��?�81N�Kf��ݱ��4L�&� ?:�5t�Q�>W@r5�BM���h��S��'�['�b�;h䅆툔a����KzeU�̭�_��D9$5*��u��N�3��nL]!���f-j?�ɄY!�^�t�=����!x��~��N�i���hb�a�r�Ɔ�[B�qN������&#��>C��X ,��,��''ʟ<��I��\���������߁�X�:u�Dr[9�x��8���O���~��T��G��g��E��Q� ?׫�%)�4t��&,��J_�t�lEj�����i�9�3޶�¶��� ���Wk��|��6��'O�+�$�`�\%��� �:���4�1�(3��*%�`6i�V���8+�ѾK=�y=%�4i�iy��tRf�"2OK���ĳu%E�^��7.�����*�OV.z_�+�c�jH	��J�+����$�ȅ�m�_>C��m)�I!QU�eg.=����Vh�ݿ_�2�
X�%½"�b%�P�1�?���^��/>��4o'-k�{0����:��J7��"��n��p��,.�Ҿp:�&��*uC��Գiw>Џ�h�h'��T�d�Yc"�����QA�s!<�a��u��(�U�`�`»W��D��}:;{�1�J�5R�Q�I�c��TR�4���A�o������o�� ��lB�����x���f8^�M��r�g
2�Lܭ����LM�|?�.�g�@-{�qsb�1��u3�%zvZ">���t����SAW�'���n?ݚE_y,��)���g�x���^R�Y>�����}���b�W���%Q"7�������V�V�{�MT�#eE���:��ր����o�ς�d�=��ۜ+�ѻ�Ab/>��nJ��}z��75 ��}��ِy�x˂�Bqs����?K!1�|��>��б�`��2��$+��(ʧ/��Dk��
�gT��K��ZX���W[�Ic�ϯ/'ť�!�g*������7i��Z��:��@��r\�������*�'>,$�+\�c%�]��鑖a�qT�8{��U�����FY��$�f�$cf��BM^�u��r��B.�}�`UO��E\�<������%� l*��eT��{�/�U.�Iх./�l�[g1���w�6�t/���i��ͽ�q |����=P��=M�s�Z����t8!V�kW=��9}x;ΰ����E�4 =�G)��6`,�T'�9BS��5�x:�(s��oZ-�/R��f=�	����m�:��O��N,'֦����g[�K6ۘp�{g����XU�L��R4GF�	߫�_��&��:���+�d�K�o�~�ه�5|뉺����8�v<�4%1K��-���;a��f(=ᑑn(_r݋����/��})�w�d�J�y�k���^xgIMɪuKx��+8����Bʏ1Q�#�$#��6���O�L�����������ܧ�\��G���$�E��k2�?���Me�/8�����<hb��=�T4���Xs0�X���s}��zF;��]�Ӌx��1Uɏ�y�Ό�$�/��w]Mf����Yo�"�X`�}��-5�i��"w[��z�X�	x!���d�Y�<�i��e;�l/x�38���/9q�qS�y�7_���X7�S���qx���(n�������剎����ⷉ'��;���lns�����]/�DI1���ҍT��	�o
YI��c�؀�����=����1���*�������t�v�[���3X'?���OlJ���2Aj��e��ߗR���Ս瓕"�y T�T�@搸KgBY�qr36�<M�)��(Wå�ޓg�:�	��RY8�ת�jd�G-L��w5��d{�WS���Vd�v{���a'<	�#�Ș ���]Z	����~ъܐ�n�Wl���m[�;�4>�b����;j�6�{r�?��o��|=�<\�ߵ������~T�0Y�"�>��J~���RX���f���| �����[j�S�`k��ݝ&c�s�֜�eIi��_mv���9rrWW�9^p���?�,!����y��
A���e)�-��5)���zn���<�����Ԇ2����f�p�3G���1}�Ḋ���7���j�i�g��~H�C^ 5���[BCml�2��t��[z"���T�ۄ_lH���B��rG���.��)��3��S&Q���<��X�!���=C������je�4	�ׯ�=i����w,D�bX���8�bO��\�^��c�Hq�>�b��l���g���Y�6����Q	`��k������D+97/H۩֟�|#�=��G�yҳ��� kǊ羬�3럆��ʁ�M����i��1���%���&$^��<�^��N����݋����b�G%>�ֶ�{BC�e`��Q;%��p&�4F�h��"]M�9�sw��˦ ���C1�
K���I��ι��ߍ�{��N���5kQ�n�)�<Լ�ќ��Dr75F!CU��_����e�y˩�B#n��� u]T�yo�]Ђ'gF̴�ia�S���]����vY�h�V�.O��z{�g�;{Ӫr���h䷺	sXZ#q��p=_V�כK����&�Gf`����t��"+�9�U����=�ѵtρ��.������=�Y]vn����Ã��L;�f�p�ڋ����d��p�x?�x��~��R���R�t��'�N�r"�rF������2Y�֮�@�)���[�E���K����ZF�U���Ɇ�A�&��Bg�n�H�wFv�7��߸6,���1th����~��蝶TEe6����t��i}�W��l6��mq/�C/��G F� N#�gq�"'���8>_K�d����WSW�C�P��������fF_�������X�k��B/?�ԇl�IL��D&�۪ %���#{�.s��xN�Lt��N��F�0硙zD"eN��C\O�e�߁�Y�^O�����zlXLW~���h>�R��� ͩ��Ҧ��~��0�/�`X7C
���4C��w�z�*fV��ۅ���N&��L����^�sS�1�z?�T�H'C������	��߇��f��&�H0�9`GK:sz��2���8OtYg�0*{�
�1U^u��	�|��Z�Qx������Q�W����ێp��>q���ɶ�RI�Cӝ\����4x���6um������d"�9ݴ,��r1]��Rq�䥍�@W�A���DJ=,���V%][M��-~���s���S��͛���lrXuha�$�eӹDrъh
��d�T��&��c���������>6�bO�����0mqw�vI�ۍ_5T.���j̿��Hu��k{!���s�����xM�������R'ݫ	��G�d�u��7F��2!R��Cp��p��H��ﳇ�;��$g�4n��l{�-OO�l���y9���=hZe�=��r`�SK5X�o&ؔ��&� ԨԼ�M����(��%���!B��_�cJMˆh�Z��u�����!WB��� ��櫦�2P�_N7�����N</��a������n�%��pB��_|p�U�,���A�w͖�o�֗fi{c�MW�Y�}�?�&]�);ILrY>q��D�O0�`�R$�iG_��lT�A��*�(��M�Y�\נ�G���.���%��B©��������� �H�7:{�.	1��߇��LoF��ө���az¡��~�<��U���O{����uyK��W����.A5��"��>[M�y1�\j��s3����]���7��@�_gZ�	Pp�0T�ŏ6M����R���%�ԍ���C~�]=\�bE<�n����b���3�;[�RT��_�^���� �h�CB�p�ۭ�F�s���n�C�!gI�1�r���d���څVV�M���"j6�����3�9ƹj|����Asߡy��Bƾ®,�T.� � ���t���2���!2����sq�4Av���]b�9B����:Ȣ{2�i9� �Y�M�k򞳪�H���Y_>�w��7���-��*�5�0^��u����Bm�����W'�mAFM�����$���U�i�߭]}*���Ma@ �SӵM�/�~ь��e�f��%I(���b�m2�)cdf���<�y���l��I��z�򈼓�9���0G�a�f뉄��L��(����+9?�M�^Y���oԎ\�������oGE.�q��N�e���7y2SP�J��Ƙ��H��X�!�åVl�0��_����Dr\�����e����f�D�TAq����E�Q�,��֯��c6�j���'Л<ŀ�g G�p1�Ck�qn=n���7�;��Ȗ���wGY�8ν��+��MI�/:@;mT!o�~7�p��y������r��Λ�4mfՠ�=^�%��� Ö�;�,���SY��$od5\+06�3�����x���n��<�')�u���ߞ�:8L���ֻ@k�/��idx��b�	�m�L8�k�8�+�r�X7�^�e��קu^�/�Ϭ��L����m~طoگf��@Ĩ�ˡ�92�����nV�],Ԩ%�:�>��4 ;��q��XY7'�H&�8�_�F������37�^vȜ=�Ĺ�����g���L�Z��QY:���k�����j��\E{56A���7 �xy�L�޽�w�phrҮe���2!B&�e�J�>�h�^��)<E�(�\�̌��f3��vl䪑��T��^�V{���
fD��#\����矬��i *��5=�k{�'��P�vt��(�07�s/��ohM�u�a���7c�׹�{�ɼ�m�V�9�ҽ��aasA���P��m�QM�0O:se ��*�8�2�RQ˩Ċ.a�|�ɆD���g�Z�q�4fæ��g?�C��e�J�� �Е7cr�f��re�7�,�|.����[�����r)U�V}FM�6_�����ڬ	��Q�f�HD+�⥝#/�'���E�f���D?��	�n�T�|n��d�Z�{{�JW��|��ɔ�Z�o�"����F2��۶�g�՘|W[�����c9P�'f�,"�TCE��B��k�Ä���޿����G16�`�"z�^�Ʌ^;�s����a��#D��0�p��Lv��FEg�Xޕ>��F*G`���G�{3�b�A��)�GX�xc�V�*L0p�7j�||46������e����^ �N�1r��ڐL�v�æ&UPN&�J��+⧣߶��2]���Z�#�V�aD�ˀ��o��M{)�4{s'�Z��%w�<�5�Q��筼i#wu�y��>��y6�W�������/�J%�/O��*kj8惠B����`졃
Y�l��d as�� �B蔚_���&1����|�$ �X� C͘��w 6i��i^`�ֱ-`Ji��sv�8Ȁ|['��(�?��;��zqd���H������/fI�2k/��ɷk��M^qF��o�ԡ'J6_��b�������9x�n�c��ww�֤i�'��:[&�x��ѭ祫0-��T�&��@�B�f�y!�ż���ژ-m�nA��>7���D���e��e���c�x�7�؀H��$W�$fpI��*��s!uPc�̢�m�j�J/���e*�������@0�ԻC����`!����D�?�-a���Zhs5=�O�O����[��4)zRDF6\��hi�ϝ��R�У��ce��cIQM)��M�`ϭ�Z|zd�,�J8�Lw��F������@ ׀ڴ�Er�ٛ�Ph�A5VԶ�z�A
bk�O><�M�\����^��8�;W�K^���1�v ��U�v���J/�oze>^�ķҵ�?k�Io��-w�Y՟7�o�����XX���ɝ�i�[�V�ɫ
6������s-���4r�b$~�:;\�MEK'"�3�j?3��3+��|2%��/w�8�C(�#L�I8o�s-�}f2�z��1=UI��n�:T�8�OÉ~�M��]���%�\�^y�����8��\|@$`�<{."/����V�do#J!�����M�^u#AÖ ��$���݁O=���,T��Y��dK�1�� �0yS����0�yG�Iמ���[��J\��+�4*�L���e;["���(��ڣ�W?J�	�\�Q2k�Tp����q�szH�y�����0�߱iHy.��Wt�t�<L����De`j��s����a6�G9f"7��L�v<n���y�Bڛ�8E�M���'�~UD����b��!Z��Ն��ո_ݛ�\�#P�7�)��'}�el_2�.q.3����e�=����&ᖑ��"y!���#ݔ�oֳ�VH��v�[�f^���Ӯ���Z@0s8]x�d�I2-�u��I�&�����:]�w�G�x�4�`f#��*�[X5�ϝ*�w �}�w�1���'���!�E���y�����T���Ų~�q*l0%�.�pŗA�ւyE!��l�w��WV𩬐�k����l�)F&�9�7����r��LUU��,3t��N��);zp�	&��*(�,U`��!i�����Y`z�1�0��6�p%Dp�|葭e�k8�zS�F�=d�%���Q�,��I�BV�2��M����i2���M��18\3�����=��vL�.R���̪�h
�"OHG�6@0� .��s��=~�A���{_"#oS�ҡ?����ʨ�}O$��4)��r�+ U,�rNcD�W���+�*��ӡ�{�;��;�-�=��8�yW�)�.�/'y�u)����_ג4�2��	=,�͡v+���	�ٛq���3��	oq�[RB�&l�U���#o��Rt\�v9�0yޭ<��`�@d�����ͦ�8x b�����k ��D��r� �)Ò%t6���l}�����ߢ�����a�B���
��=G"r�Qv/rɄ�?�T�-���Ba�%mi�k`�i.�9�wv�z^�h�F���(L,6Ȼ��:���D�Q^9c9�x6	t+��v�ʉ�W��:�!/)��K����F6�*W؇ �+�������q�F��Eڡ�.����k?�<�_��+����h��"ϧ�"!�J�,C.(���νD��0��c>،qؓg4�ڣ�`�D*Jl���#uue�(~��4��N�~<�fz�'�N������冴GgQ)��Y���H�^��]A���@����Z�s2����:�����\�t,�˟Pu�ZFudSP�6�3�X`����b��z��g|�( >�ߠ�p�S熟�i�a�
ı�ך��i}�/͉?�R��j n��BK��|މ�K��2�M7~�G�Gy��;>6y9�!N���+��q��&��jp��7'@i��@�Ázr<Sfv/'��qV����=�D�R��E�}p�f�:�!��z-$�E	ZK��<-�9ij[�j�~�]Y#��m/�mZ����
{�%%S,��:�O"�O�d�r<aNWf��.ۻw1����TQ���"e�����gl%��3[eݢИ����K�	V�T��r%��I7ݖ7&��Pj_�3|:�rKF�N6��w������ W�XؓQ��{Ew��L"5�W�����4��*�/���:���ڙ>"5`�+��:u�k$-G	S���sn���	a�>:G�;�� ��U���3�$V�I,ꈐ��`�|��-�A5�a��Y� ���!���1[	��3����Kbj8H>	��cU�a�;m��h���aD��]x��4/67�VH\�3R� vC��Y���2���k��uC��Ϥi�.�j�٪��-���{��U
�HW̯s?T���L���z���<ٝ~�^?����T3���F��H��?x�n��#��Lm��mx#���1R���:�f��%\oQ)��JlƝ�7l�,*)�_弊*��3 ���z�:p��������{�o�P�q%(�/�P��Ҡ�dr7gB��\'oZդ�\<�c�z0S8]loA��W���T�N}��o-�^Y���[�ã�^�5	2�3ZC}���}�����.�	9�Jչ��Dze���A٢�Z<7
��_�R�ϐ�v��B-\���QVvL̽)�-���$D	D�,�`��U尘gi�$��
L���_`�,��
'�x�2�di�e�������46u/���N6s] ]_�HU?�	L���<7�{%���d��?���4�:5j������q�^r"�KN��PAݤC*�Z&_l��9���%K���x� RR � d+r��s�+��T"�m|����׃r�B$>���B�J{?�f��9��f��k�([p�#j�'��7�)P�q�޴� I,F B6��ex�����F8��13��פ�\��]����U@E�>��[@Ji�nP��.��A��D����\�c�󻋿�w�G<���y�y�y�wGر�݋�_�?���Y;���`I�T��=��#�����6[�>�yhv{Ȼ2�5��G �5���5˪�'�+��-C\�`iI}�	�i�z�7[uA�t,���D�Ju!���ъ�������H�yҒ��t��*?��:@[ =\Z �j1��0�n�}vӜ3����_�qcoBlR�!{�QaE����E�j��=\D���~G�aP[{���Ta�:~ܲ=�Wf�ӳ�5?Q��2URW+X^TJP�"��p;7Py��YQK]���n�$z��G>bu�h�ۉ�E� q��@�����N�n����֏4�ی��
�*])Ӟ
�Fi����v}z�Q�}y������)Sn7WVS�_��ō?k&�ҋ"t�ݨ�M�p80�X��$L�O��A�_õ�P�R)a�1�ʛ���9�&��D����'o�"@}zN<��[����֞�-�~?�]D�����B�{���?X��{v|.-4���hnX���X��_��]
^������Vc���G͖��󚚤9]�c���Ρ�$ߞ��8؍�.�m�Is	���t��s�V��s���cd�,̗�rG���.q~ b���ym)�υ�I+Hq�������ϸ�H&�fj�ʐ��
��I��ɀ+�^��;�*���D`S��1�ƥ�N�G�r0���A ���Ŧc���H�Q�4]$�џ丟�s[��m7
)6
=(���u}]n���S�oI�(����Ȩ���.OR��׳N:pձAg��CdoE���eͻ�YR�S��u�b5�ߴ;����NM�����U"����`O3�:�m�x���#�Ys��c��VM��`�|���.7z!#;��̤ǂ�׈�������Y
�l9�����N?�5k �%��(l68K��P~�&s�Q�3�&PP%T`�`��f��T��U�cI���Qb" kf���LSe��W����E$������o�Tv2������n�'�;~B�6�M���%�Ǖ�;z����ܹs��6�A�`��C��)��>`���=�}���Tι�}�D��qB#��ۼ'Z>��F.^a�:2P�V��ݑJ��W�s�^{c�d7�&�+%l�{�"��z-MLd#9+�P1���"G��)��>����J���7/?��@r"�q��f�T6q3�ݳ֔_���p�*�Ň�>�?l�W��۠���Rއ܅Z<\ ��' }>3��}��[�D�5U+��kQ~��f�J��d��WA��`�[�.��`O0�	��j�j�g��s��)�y(o@L�*Zw���E����,�Tgu~���
ے�1߹��&�N�-ov���f��\��"G��nSC,�ր��ki��>��I���3����'�H���X ��f1u�;�4����Ŭ���~���a:=��xOB�nN]Y)�d�<�@�Se\Xa��6ﯖ���륏g��	XT�hēK��Pm�Do�ԋJ'B��9�;L���9�SŒ�IL�p!��l��Q�DK���_w�S�G�qػ(w��Ү�����R�_wr�U�S�I
A�ِ��p�RuT>;�
����+����Qˋ�o��M�Ο����=P`9�咷��_r��P�W`ć�E�`��ǫf*��vCr}�/�� ��(�=
b�>�Z�3�zAx9��iw�B��&��s������
u�P�Z5g�l3Ao
"��Ɗ��Q+}d�k���D�5 F:��睳=Rp�|E|'��^ڊ59^aY�d��<��q�����Q?/F9͸�3c;������?���|�n�
ZE�/��o[�(lM�*�n����S�z�Ve�0�ɸ��S/�(|%�WF�;�DS�En��!����V���t�5�ϙ�g=a� 7'�x"c:�&9�m���%~��~Kp�R�*�Sܣ���;%��Z#A�xCe2;���wӡ������5�?w�h��*�ׇ�l;�ۣ����m��{����Z��V۰{�0-����(�%]�g�����ͳR���aPݰ�1�%�w��DT?��.������tY�ٸ�+��]��m���+ʮK�O���6�����J��S�ӘL(������}=)�;#���6C:V4!�"�y��q�K�-�4��ƴ���Q�����?(�{�l�nwtI��&��oj(GS�	*�a2�hհ�HB���-n ;|l��ޱa$A�ئ}�	,Xͨs���b�� ��q�q�(���QoX�<R�wk��o�@�nu�zῸ�~�%�﷌SVS ��km��!���J�1��1�k/�������P�3���[��Q�r ʲv�%�a�R8��7:Ȼ./�c)i�4{�y��W�ʞT��[SU��y�!��g������x��ٟ�:I������"^�?�����M�eP��2�!j{�K%4�lv@�B�[�@o3�J�t;����H.3�;�f��9�~Q_�����k�ť,��L��K�Z�WF��Z��b8�l17#$�R��/'���y�a !L��w�eCQv���Y ��O���T��Wx��y�u�����y,��L� S7_YJw�ByH�캖��Q���nMY�N�/�%��T�xo�ɑ���O�h�d_e����_�$ ]���=OΊ:�m&�`����&!���vY��� �#��'���S*<az�w�J���^���Җ ��T��H�Ӝ�3�_I�'<�P�[����a����O4�!��Fm`���K
\��R�3���n�^zR�&K���|��+媎c�2���
Ȟ�j��khI:�1��rT�5E�>h�u�v����|]��JMp��ν$�����������\
�*(?5{)&Me� �[�w�	΄�5��:x��������U�I��ن�hק�1�Vm��57�Ⱦ���d�[�m�?��*Nϩ��W(L�
�� 
�$���Eb�4o&�\�^���f;w���nӁ�7s�I�l ��5�����zQں"��5jX}zݫ�K�����at��T�=޵y������������m�*c˼�Y���^�rWwDo�M��`��T�k�l���ˋ{�a�
nam��u�WX�.r��5;�8�.fgD���.�A��� �̈́����	5��FO4 �X}I-����D`v@��x6S<mVw_��ց=�#�B �̓[@a�H��D�j��,;G��!�DWhY%���2�D��C)KV�����QX��Ϡ�{�6M�#ЪS�r#}�5e�]���̳�>��\PIg��q�w�������%�#@Ȅ&1��K6���fyw�< j�#R4�MwE{���;+y|0��0��U���d�R`B{̸5X�/W�x�4s�!�ީ�1�Wr����	?uȚ�C���]�A����;y��x�Æ光��΋���w Cb��uM;��0�컮�\P����#��̥|�r���I�,�M����op�6u矡���Ԝ)��+h.��/���l �w�g���s�H%� ��p�S�>��2�������h�m����I��`j�a�qo����O�y6�I
���ￅ\����rh �&mo���m[˴��:��D�TPc]�fu�]��&7����$s4~H��� �3�x����b��Y|�d��0�ZB������$s��j��]��ؽ@��
W���`+'� �򛻊_Y(	��D�2]��*f��t����Ӗ��ߧ�cM�~���Tɯ�Ca�X�R���r^3ﭫ>�2e����*GU=���t�++�v�_������Q�ռ�Ű�ϏА�W�Kf4mh�Sm��kD�/��,7>=�6�s]�q��
���TS��Ǟ�ŉ��|�T4A�̊7�F����������-�4�}�<��V�}���{%ۨ����wŗ�ַ_~{��䈠���o~�s�+�]���Ex��jx�'9Ǭ��u�9E�#K h2�D}!J���G.ʋ�#/Z,�H�g��6��o��x�M��$f'�P_�'y�ߏ��?f��)g�/V�v��qw@i��dqϪ��ßZ,�&�t;�]w�sG��[c?������,��㖾N&(�+��iv]��S���,"� ����yt�T��5+q�0�ǭ��0�<���w��_|�G��y����|�e�@�x�R�5��a�b���J���±��=	����	�*4�	���� �į	i���ws��O�$HY󺕅,���p�X��C`C�ZB+>�{pY�²�>E�ڒ�+��/xv0�Ċ
�{[��:�7���r�����SI�O�Sr>=X�s�����}����2xT��$��D��:�U�1jI�������?��EѹI��C`tAO3R:�Y���4����B.��	��@&"��f]��>�ڞ�0��W p�}c��J8�m���C���s����⍇���<�H�?sch�}	V =���`h4�Q�UD[i񓿖���^�r��Dk��Y�/wϧi5W�te�n��)�X��.!2I�UjW~癸f��<�g���hA�CS�l�\�=��i��m�ӟl�{�oG�P�9檁��P,�z��&_n�}�㗴��<-�m��ۂ�D�	�=���������~���T�����6�/�J@?���h7���xƞP:��5�¶V2\�k�_�C�~a������Et�!@�cdUm
�[�<�%��^6[�����lq}�BbA�˿���j�̭G��I$�h0@��g
t�d������M��W7߬-�߳ܵ�aP�pT�k�:}0Ud(m�Աt(�k1���/�������wx�4m	s���x���Ҵ���x(.�
���Rg5D@%�d0%3*a�Vr >B�$ ����h�_�S�s����Y��ᵷ�a�N��U��}��ѩ※�������(tw��#t�aJ�?t�\��d	�{��x�L@o.V��׺��@撮��c����I�L���nh0����^�GD�O���J7fb��,�o��,/�
��b��!��?u+o[�П��*܅�!N��:�0s�B^��$�X�}�s���\�0N#@X�W@�Jy]�r�A[�i����E�Cm�����������Ic�F?��I-ۓf"p�S�0$wg1i�6��/��k.��%	qm�w\J���ҵ��v��yZ��=p�~�k��l�6�le����g�U�n�u����O����A�G?��^'ig�<�g24���~�D��5:��s��Đ��ؙcT��r�����LM۶���fןe4[xHE���N;�j�����B���|�O��'Hw��:R������q\������P�!�<s�ω���-��H+1��=���*7,�A �%�7�/��H|0�]��>�b��Ex_/Â�9�C�r���݁����y�d��9^��8�����O�M#a�r����W�w�T��%�=����Ć"K��zō�l�ڑ�P� =����� #�l�	!\��C�F��)�j�ޖ$Ⱥ��>���=�ј�ܯ_eq%[����f����C�"</s�/c�Yx�]b�^ R��g��*�wl���V
ѓ�<�UET[��aZ��9��:]����$9r�j8ѹ�R�H���Lf���H��$��� ��r�� ~�=����3긕�&^~��F�����M�Y��WЃ��r��6�t3��͚�Vf}TNoO�I���������sq������0=�F����zm�|��z�Ɨ��>Uˆ�١�m�fO�yC��ǰn��4sg�Ƭ�|���eh|5���nA���~����i�u%׷�lAL�����n{�T�*>f����]�D�rG켤~@��o>��z�"J�Z�}{�h��[Wg@��\$�:����5|4�y��Z��i�>[�W�G%�M������CMjؠ+2=l�ea���_���SԨ�[o�>�Q��/���s���_`Ӝ�`.��7�o�����"��s�V�B�F�sx��,a�T�%�L��?�4p��$���o�S�?T�7�g*kq,P_@j��$Ud\�n��gy���㒔Kd�Ȱ���Pae�4�}i��#�Sd�'��%�\�8�����H���t��ڹ)�D�a����vν�����������_���$�������C��ta�
����K$��`����{3e�¹j�N��$d� ���m�(�k��CD�`�E��C|�﷋�s�]���S?A��������-\�Ǭ���ݝ��?B��� O}�	H,�y
q�W������X����9�<9`dvh��{��z��I(��șeok1��	I�pT@�gu�q1$1`��nQ����`�<�H�o�A�z�|�B'��K�ɳ& M�[ض���g|��9 -{2l�/]���}+¸q�P?�}��_������� ��.qi�4v%��w"?�����D�e����,�}��~�^�~6E�)b�?4d�C�g�{T2'
���+|�{�}LV���'葾��!٧�,2��"I��m�P�A���n0_��F�����Ud�.�`���3N��e{q���S@q�j��o�w�o5���g}5C��Sl��ǃ���nV8�G��V��+ءx��T���5�_|�H+o���1A
����F�	Cg�P�씿������ً7`e:"��<������~�ㆥK�($����nΰ+�M�W8B���G�y�J�;u2�~::7�UM����o�vĩ9ˆ�xgdiA�s��q���D����F�	W�FSA�����M��I{���g�Ұe���{���w;�&�IZy��Uv"�Cϡur�9!e�+Ү���ŋI-m9��}^�%'�Yن����ѾSU�p�&��]�)ǵ����Y�|��ma�s�+��b�\�k�)za��R�]N�hP�2�k�r�@(e������a���B��Ǿ��w~NsF���y��*z�-�.��ـ@��ck5y3����̶b����Ә}	��������#��}3]u���ֆ4�w��tSWp��(�ν�*=3q��{�����-��}���h8K��70#p��8����V�m7�6��-9��3&�ʥ��i���>K�Eqh�W�]6��)�x#�hE�Z9IL�^XA^� �n,>X���!���'hW����5��N,��A�c5�����Hd�Tta��/Q�#�3g�J���� �
M2�\c� m}*��֗��i<ô*���I8�@]~V�W躵���캺��Զ�'l󫼨��{���t�����N㋿�Y�Z�xa�fTԜW��/帺�#D@@�!��K���ki�z��F3�-'2ܑ��'r���4�
��'Z�I�<9D����"��l'��!@��u�ր�E5�zi�q��s�k�qȳ����);��B
P���%���z*�7�{<#:9�~Q?��	Fg�å<���xLZQ�
6�qdoU��v4�P���o��	F\TQ_d��Y�_�V�}Q;M^uf��Ӹ������7��;�eq���+���s���G�.,s��ޝ6'����LS�@��kM����R�&�$���ר���@PN>>�%�0��A��,��F� EE�JE�y]��BiM�O�2������G�<ά`�	�����'��?,]�8���t�+��"HoW�pA�Tvj9�}7�x�?-N,ˡU��| �LN���tX@r��R�ɟ��2?S��Xۍ����ͩ�ޔ]�C��p�����Q�A��%���h�G�c���@���3�#������r��)���0��'Q��H<�7䬄}�8w����G�<9��Ǒ<y����`S0��0N;�PT�K��c��A{�#V�HZ�������I)ք;b���� �|b�����d*{��d�B������,=������ۡ�7���<��"A��>��4�my���m��[�˕ \+
�\)Y�ua�- I�q�,?q�M��.�K�j3��������^�f���,�>{���<ܗbı�'l8�5�EEI�ƾ-���$ŗR��Og2WBmWIMM9P~���k;؀o*0{7T�	��H���ǎ���*4�Ȅ�íFв�ܖ�T��z~���k�c[2<��c��b������|6Ԑ�lK�4>�nM�h��:I����^��>-j���v��i�������1����:��دW6c	���L.�k�͔�S=���0Xq�W	:������]t-g[�#Ϲk| ��V�G����}ݛis��W�������׶V"���2��Ϝ��LuQ:�Sr5��)�L6VE�T���#0k�兇X6xh�k ��oO͗%�U��~�jI�'�i���l�<�[��b�rc���9��������w��Ȟ����3:���y[�(�xl�0��+�l:s�]\�� }/���4Jt6�Bƫ
ו����,k��!2߃��F��K��i�m�^�5�&�V�+@�C,k�	�-D�/�����!j�g-�5֨������^tq/CtG�������dH|��Fb�$�"������n�H�J��S ��P�Q����T#����)��T�_��V=M- um=S$���>H(��ê}�|��`|��ā���.ԽC]�&,��A�qM�(g��O5B������[�p�Z�!2��t�����d�������<Ej>����P��4d����6���<�y�ۑ��k}��>ր}w�1;ή��kt�r���c{�*iD���%B�׹!��@l_ΐxo��
��`��j�*rУF�.���o�) }������g#���!a����6E2�*�TL�Q&���(�W��֌��*dof�'���_}�D�ٌ��%�,B�7���h���k#��#7�$K��A}'l�J�R�d�rkY�����~��mZ5td9��rjӷVa'w���+bKi��a��Y+�9\��o7������
���h}ҕ��_���]ݿs���)o{E5�bGF�c&<����=��T�:���rFg��������Y$�=�@��E�K �$ҥ�T�J}u�ܘ亱�O�&=W��ǲ|��d����o5E�\}�/���L]�?�SQy5�^;�\�)lj����+�J�+�%�W��X���R
�t���$��ɤ�/�2E@wNv�z2ֽ	2H��a��IQ!0��wc�DT��Q4b�7jrhp�^1#���V�q ��x��I�tG��E	w<�&Sd�ov.�ayp�jrSyF��@�+dx)�Z�4c��,p�,i�+4a�?�;y����<�?��+xz�BO����l�
�z����MYR g�s����*�7��^�����~���O��c�ޛ��	��	_�0��tP����C���<�g>���#�oy�zrC�?g�\q%�ms;�T�Ga�*�f/_~�S48�e�������o��#�t m>@Nx@/~х E����<����D�m �T�c.ZTE=)h$h�Ĺ,?5ΰ|�a�Zr�{��k�EIG;4��Oʈ�N�B`ʺ}�����Wq���;Ǟ��w�eIf_L�[�ҡl�a�.SJ�d�������\qe����Ѥ��l��2>,w��"]�S���p�T��t��X�F��z\B8��~xbx��7MI~=���2):��=#j�uQv�ڌu�d<?
n!I(������P��j��ɛ�2+_\��~����툝��A\N�]��!�Y�
ƻ���� ���H����-�x����q,ya�(=�Z0�1���[���".�7���wfyzaj��q$t��@��cِ������u��o��� ��s���F�#L��wӵd̪B��W�o�@��{�P�3�� �'��x���䱽rQB{�m[k\��ʜP��4��࡝�V�Ե��X2Zf�1�R�D�!^�
��e�^]VϪ�X����Cy����������q��������D�-�Dh�Hp�Nt5�m3f�(�NGA�@!>�_h(�޹��螎���(�4T���z��G&�+�A�)�sI�܎��yot�*#+ǁ��&�2=���sS)����=�`���'Ǡ��[�_�#΂�hAs�xﾓ��L�o��2�@b啧��<�x*ԓ\D�Q��ȫ���~�T�p
������g���X�����X2H�����͜;�[��l��\�t:F�o�8��M�]K	^g���)#�� 9�����W���г���C�OP��~���Z2A?\N�/�@� )�����#�GX-�{`Sq�[K��K��VK
�Gy*��'V8�������4��*P���� ����xXq��{��%13^,<��)otHo�m����u��/ĪV�ցa?V64����e�	WR?o|b|fs���E��������fd-2� z�9��p�t�[����Rϯ�����h�,s6s�JC��,��=��*����	�i-�3�䮗���=��8L���Oջ ���餑5,�H*��B����y$m��U���^���@aڤ^�휐�(=O����ĭ��Ӌ�ʋ�k�t����*�w��~x�8˙vs�I�x��}��z:Αz��4F�p�8������B��P|����,-�Md�ǐ�c42�>F���8�7L�9�M��Ĥ����1�������/Z>�{��*���	�X��Z-�֗��y�#ky�;����1�)�|U�L%�*
��b�Y.���֫�u� �ͭ�o�����H�W�"�/.����	�oG��R���Dl0��0��t�-���& ����f~����f�z�)>[}�����R$bׅ`�w�y2�l`�M�b�G_��A�g�I<7��n[p��?���[���&�:�6?�~��C����!{��<��G�E�b��Ix��P�������E�?����܂��u'���w˕m��t �dT��w���|�k�|ߚa#�tA:�1�X0�����n�6?��)3$��o��k�`qn%�/�y�&��-�h��y��v�ܲ�c̦O����=�zK�3�t�U� \"ha����P(�"n�H`i�z	?�}Fq����Ф.�����y�����D��љ,V�j2(��u��ԙ��zg.���;�P"�n�ac�5�ܯp�:ŷ|o�V��ai�A2�@�S�V��L��4ih�"z-�M��� \���`�~&�q L'��n"���q,��������l81�NK[�%��Q�0D����p����`����R��w�\�A|)���wԱ���©K���i�լ���مW1�>$u���m*L�������YH�J��&OFs�v&��r��	��8	��)��T�܌�N�&D��	+���{�H�/<��Y�B`���xZ�n�-������;�S@�qy��f��߸{�7ҥ������_�U��ڲ��иm�39P���"[��@%A
�G7�����1�ͮ�ݺ�uW��0 1�?�O��|Y�����V�'��[q�;�|���QZ�t���;��w%��ϝW��$����e�Q�̱��$�Ϩ�������B�𷗖�=V��?�`�<*;����>��.�FK�`��s���o(��~jK�σZ����	���re +S}��UAуn���%� ���ĥN� �(�)�<A! 8�"�q��2���'����Bk���;"���fZO�*��.�LC�Y[����)�>/���r�C�]̆V0�:9��]���d�<��l� ��Q8�j�,��v�f����9��t�^��&�Ʃ���C��V<x*�y Ρ ��;V����Z䞧�W��s�����4���;ɇ�e�&�}Po����~��=�?��7�F��F�� V����@@L��]M�kF ��{2뾸\��o�L�j��f���UM����EKL��ޘ�
A�x�Si��y���9=��B���� ϑ
�e)���Wjj3��(��b��۷`�����
�	j�@'zzz$���wՒKU�'b��(7���N�"�4�L�4�!kj��kM~k�Wo7,ede-�yK�4߮`jR��������`D��lEl�ɶ��m_��Y~�o'�&�$�\���������k����B���M,��J�q�o��u�<��V�_9{�a*��d����3��!�9;�J��wB��\ W>���=+�DC���W����h	l���w��;rBo�C&d�?n�v���g���<͖�5���$�1G�����*�f�������?�"���<[��`�\:���K�Ig�s�Ԅyn����Ț\ �JZi�S'�Z��6d�n�@}��+��]�I�Nc g�+�:T[v':4��EU$����zV �h�2��	�N}�*�U���j'��C�\с��n�h�k�{Pa2O��7u'6��4�K�U�\K��qc���#����CʓFZ��?��O~�������H�o�k,B��ߍ
��D7���p�L�Zx���#��DLxar~9r�\�״cEG�)���bC<�&��ږ��zz¿&�i}��d̎�>_�G�TS��lwm���`��Z�{�[v��?�Fv�|-X}�CwqH�)%������?�:�KD7����K5��]�`�7�����<n�J,(Ŏ�K���g濻�(癩��+<�B*ž��J�#��C��!�5I�'��X�,R���j�K�\�4K�4K9 �.B�h%�7oB$+��F��U���h�㮰��V�� �b�9T�����L�3����Em9���$�&s'ދ(.�o���ȸ��U+��yU[{Z`|b�NR����,AUT�!S��P �1�E3��tOS�7pa:9=I�~5g_�e��&���������`�Ssj��t|��7HЋ����έ��"��Y�k�gV>5��㭕Yj�x�����srg�����F)A�5�W1�������n����:�ඟ2�U�*�g�ݤ��,�]�s������;K���0=���1R�>�+�<﹊��7w'�NN�,8�����`8�R���O@0�[�C���ֳ��K����5��Vh��߈w���ڟ�nw��n�^�S���TV1���;�d@���ݣ&DY2�u���:���Y:����o�����u		L'~�੥�k0�*���
U�Fu���i��R�Ξq>�O�MQ��/L��&!#� p�G�l��r�šs��J�G��b�;��
�wz��|er/%����Dm��y��Y �OSS��.��4������	"�`��8Ա��n�]� g��p�?�4�6�����I:��T���xӥ�&ߪ1�y�"."7@=�B(�N�+�0�ӌi�ge�Ҁ=ȁ�W�k7�����cLT��~\�-����⏈+�k��V�c�,���!�����X�U�$~�_Xj������
5��[�{�c�����Qk7��8����E"8��A1JKBA�s��uwC�M]0����1�%�!e�)���<8���o�\�� @��el���D1+���!���z��F�`y�`Ps�FPas3KQw�̸�f�ݞ���s3.���/� ��vv�Ǧ���L`G�t���m{ĄHT:��df����fk��ؽ��g\�ӗ�1�v�v������q�S\����L�-�Q�p�w�a!���_�����>����J����P�s�F<Q�r�I���xs�:�m��?1
�z�~%������r.�l�����3��-w��K74�Kҫv$ȹ+�
ͯ�h��Ĉ��CЪ��)��(���h%V%k'M�4	���������<L,O}W��,�r���ܗ�j ���7d��w
��N���
�6���$�7�A i�w#7f�`��K!A߇��f��~�דXW}u����d_�������S�x,ȵA�V=��F�W��^f��]r���$�r�KMx�2��𕧬�t+]'hȶ���m.�r�`���.M�kN=c.B'������`p	9����P�J��%"e�<��J�R6��%TS�h�Lp�f%�����dH�z�=	:e���Q����eY���{�/]�S���K��V��~�';��~}��LCA���$���t/ދ<EdDCN aG
um������Xj�`����Oa�� �ʈ�^��B����W��f� �b*l�O
&������_D��q���N����Q8� a����)(��C
�7%`s^g:��@�?�c*��2韃�<L�&��AV��(���i0s:�^�-��ľ`��!���]�8���V�6�� t˾�%��sAO�Ȳ�f?t~��_j��<��D�9���Q=�JG@	��tr�2�c��w:7��p�觰�G�"xxf�m~`��L�{����)��PM�?S����?5xj�$���{ء?�p	R}_�v�<~�9��c��/�])0�d[�^��_���P�t?�[P�n3��f�w�#��C�P�8��Q�T%2�i��U�|�F����0����`ch5�e]����@��+����xJ�9�|컎�")`����ճyd;�-t���Y���>n��p�W'x���_���w���ʢ�*�q�P����.��A�Ƃ��|�i��ġ�͵�����T�{�_�k_�sE��"��i5�7�����(�*K��IֵmL<��͢�/��FءV�T�%?�2�D,�%+w�y�c{��[Vտ+�+/N�~/�p){�'�:�����LY�+k��k�J>�>�����H����ʍ_F���=�q[|)�G�Կ����"��L�n\�R������Z����6�����$ߡ�ש���B�3s��J:c����~zt?�g$dkaS�[/�[�}�Kq�>�q\��࿘<��U��R����_�ʐr̍Vs~1�&���ㄦk�D� �6�&t|~�Yt�E �������=���(D�A-~�73��_C���r?�<ŖB�С��g�*ǜKǹI�-@Q�D�ڈ���)��i?��T̀��<*'�fS�@��|~�jo�UD��e�9ڍy����%2��KC��R�W�@�4c�[1���!�*�`DSX���V���������J�ogv�F(S��i��$I��Y��c��Q䓷����D�e��f�/O��#F�q�-���Y- T�P���ˊ$\����R���!�����;�-���M�·a?I��^�|a�lR��yL��p
��&nl����i.,��g�k�N��#���MG���d�n0w�Ͳ7Z�G��I���\�B6��6�{ӹ§~�s�߼����7u�
����1*?�ȷ�e�`/�<�f���~��D�1S�a`]�Z]p%YB�F��GP�L���ۑpo���i�rm׾J���/�!�p��� �yi�	`NF������ej$x�L��tC߇�vN�V_��9��~V>�Vt�	�S梯�%����Ű����^�E<���Zv����EU����$����w��sʂ}��7�Qx�r �b8�Vκ�s�Ȩ���e��7VrN�8e%n�����'���P�1��ϩ=�@|d�z�x�o�G��.��� �}$�I(@�1�@�����/�\�Éb��$�l���V���U�3{���JaU��W���>�	�d{u�Ԓ>%C��m���r/��&�O�����"�	e\'َT	�����/6
�W�}�[�����e�g��0��J����מq���> ��2�Bʍ�
�$^1��W�UX�d+�4�v4�7��])�=��n����$/�o֞�v�?Vº[�
V_�T�ˬ�4jp����]�eRZ�-�cR���k�B��ja�5�����@v�]H-ηza�r2:G��\��yK��i0���޸$J�GN9��e��G>�r,B�o��9����3��9�T��FHpr��Z��C�1�-�~c�:H#;kFQ�]{�gSC�J.�l�A\5�Į�4�w�{%JBv~���u�N�ePyk�<��9.�i7���Y�ȀH�]�+-��K��;��Q�k7�6A�N�������h4�.
Kl��O�[Ǘ�8��#�.���W����=ݫ�ɂ����-:!�0��ɒ�ja\���c�T�&����2��@�>$�Tg����V��V����n������p�\����qA�bs0R��I�|�*�0٥p��E����Fa�^0�zE�}�ֹT��[Ȩ����Hw�=2�$��d��� V�">���5v���P���� ��c���FF`M'��@�[z� 2^�D/#�����F|���7[,��?lP�z��J��\W/����FK�S��Y���44~y���-���P��',A�.����h	�A�������1J���1�����i|`��V�����H=��A���/ki����_T�*�c ���}7�.w��[���E��]� �.�d$�O�{K]h��h8�����==��(����� �����,SH�|��`��n�ͨ����!A�O+^�OyE6�3��Z�*ë�}5���D|-!�*�t̸{�B����n�����Mi<#/jܴn��ot�)�8��G�gFms3	j�]���&�iR����S����/�"D�O��h�
����(LW4z��FF[p��B�ߖC�l����۲�.V��gvH���2j~g�eQ4N;����%ْ�+��+˜p���0[^ow�uNݝ��앳%4�߼!U���h�V�����/�ٔ��/P�D.aq< +��(}Z p<��y��~3�����F��C��i^�2E�k@i��%A���Ōu,Y�\l�啊�B�  �w�O�2k�`%O�U�6����?��_�Q�s�)0y�C.�&��z�@�M������N�P�h�TF.	L�HK�ŻDf�vi���������*��<���W�#��8F��M����P�D}g ���6!�.�!j��{ｋ�D�V���k�轷��GYK����X�+����_v�9�̜k�k�7t�2<R�wQ8�왠��V���d֛���}R�y������dϧ��%����k5��22X��~Zx���,�ubN�)5�Iه�}@Ey�-����L�Z��R��^���ȷ�w�q9���;���k%���iS8�����h��4�͊��*��yW8ty\>�C�9qsN#(�4U%����%O�-�C4	[9�>VʍG^w���B���-�(
��ͣI�xu�R^��(w}Z��И��B���2�%�"�<ӵ�$������Epn�k��(��b�
pm��1)-��U��nk����w�	Z�c��9���ܒgA�2�����ea�� o������RD�5�0w�a�J���(1C�e�/���'�ѝ9"���%����p�\�y��/k��s�w|��F:��4hǓ�'rq'���c���7'PF,[�Cګ,�\����=o<��\Б�?͠��I 4Usu!�W7����^��(CMqľ�0.���Q�[������O<%Gr�px]�����<�P5��L.��!�[��I_>*5�O�}!�u}�BV����]?����n�w)c|~���Y'IˬO+)��0O~����/�O<�8�a'{S�T�7�~��덩�W�m%� ���Я"
����t�	���<����E��� �6��s�n�&o󿀼Ws��fd���l�u�{a�+{窾��{BG6#�R!s��.д ./���~��N4��!D8z>뗔	+�E��Ԇ��(r�"^��7/jK+J���|*���@�Y�O��g�m����yH���h�4˚Iؤ^���F���Tt����,�*������"^A���"��?�QkGAb�Gn�������FB��MC�H����]��s�U%y%��Um��W�
>���O���'�6{�,8k2}����@�<��S�P9���L������eB��F��K��	P孈�Mg����za^藶���C��2�A��Y?���U�Zoc��8��:8# =��^ �/��g�2b���������Ž`�阴Ư���_���[69�(7�r��˪���Y��$�����;:s��6�wI�|<ُX�7gF���?�|�k΂��JU	���U�[�8w�/C�K�C+\�����ט���Ž_g��4}��BKg>�5T-|Q��7���Ȳ� ��M���>��Eow�('����#�>r�����R�~����� ƺro|�U�_�'�'�drƆ���yg�$Aav���U����3\_�g�;���o���LsB���[-�l_�F��ZD��	�ϣ�v�T��^�Z��ȼz��]��|Y�2O0�aYe+��v��E}���'ѻt�V%�g��A/��1)����
��~���ݐ҇�w�~��Rk(��+��ZR�T�ǣ��κ��_6^�I����i\��Mb����Z��G�����豧8L~�4_�~P��uV�K����nw����L󭵘��s�<uf{�����]�� X����Э��a�iF��Ҵ��-�[6���V�>9Ր�|��`'��)�Z��	�����}V��,����a�5)���Z׋"���W�\��)�=,��.�gO�!@�����i�fTMr�v+9��{(���5��!���Mf�@�)⨦R-î�,r7�%��$��:��B��J�x�pnE#�F��F���m? �n
���X�/J��� 3R�Ͻ/�v�͐2�Q'e�Jʆ|�O�Pc��
�ł��Cˇ�=�V�T�
����	�?����LW��/OF�0�y�xOTe���a�
����`�U\c���ؓ������<���v�J��pe6����mÔ�V���Z����e1ԉ��Mzp7��Q��t�'e{��_��Z�^��Ӊ{�Ŀ�À�K��p��HuQ�@�� zC��*�Bye}��B�;�I�k*K���e�W���k�M����=��
��G��6:a�5J~J��G"�W���B��{�F�fi����L@��~׺���$(��*��T�O�״��n�u��O��	��%�ߚ�W�|W{M��o�OhS���+��}���/6�<M�⾪2����!�v{�qnRn_�t �����X��:}���#��j��� 8�*/�mSN�2Mޕ��g��4���b��p���|���7��h��N(Y-���f~c�����������#�K���n},w�5�t/R��8��y��k�+l87�ﰸ�G�!.��Hj�ν=�����1S��0��ګY��0L�K�c��E����?v6��Vƺ!tY_��D3��w���$��*nL��i�P �RE��j�}.��E�i���ެ�����nf��RE��W�=L��UUy{N>� |*m��%��)z�΁,�������v�F��طU�h�8��$#Ջ�~��t��l��:���=�9�� �k�F��0�2ǒ+�a�ν۫����y�����/x 4j!J���0:��ذ�Q�!��r��'���Lӱl�k� |k�v�2���XO��|'6S�+=�̒�v˪�n�"О�~?O#- ~�_k��*Dx�@l�زb(Si(��*�O�(Gp�c��ɯ����HP��oW� �r=e _�w�@$G�(����"�;�d�T���ӻ��6	up9S{���4�]_E,쉊���l�`�)+�!�5�pF�}9:#ⴜ*eE���~P��a���jZ�����d�������̿7]��W�i�7xG�TY�5�� D����5���$�Ф(�5�^R�g�J���j�&.OQ�m�En�𙅏������F�$�/R��/�3	U�Z��'p�FL�g�z�r;���mN���ۈ�('�f��%�ڡ��Vk϶b�S��4d�)����H��=6��i��p�ȧ�.��.p�'�b����C)��Ȧ��
 �O
����0/ձ�bU��PD�i�3E��~���%K�NC|�#�YnxF���L;��`�O�ګ���Rg?�m��wTk�j(�WE�fL6��ؿ�(v��9��kDː&D����&�߱}�h��N�\��/��OX`S�"#xu��&�QN�Od�W���_ <�].i����S��Q_G���0=��>�Dlo�<�Đ2T����~�){��R
�4l#�M�_�ZPT��O��8�A�jZ���:�V��r�5X80��QK��3�Hd�����A)��?�Z=r�u��ܐ�>sO�zqO{��:�ǽUq��w��U��X����Fgk�[��i~��c/q4�iF���m5�@0�$8/ܘ�n(c~s���;�c�6×��;������$�-�P'���CA��b����_�������_�,���RƗnIs1�κ�� /JӖ=��)�Ď]��gV5�q�@�%qj���u�� ��1h�-�X�j3)��W$
Տ�@ �Y*Xӗ5Pj�Z-m����+W�{Ru��l*�շuVX���8>��ϧ��&��o���w�������v/D62=��\;ę0��<)nCN?�a�洔��� ���7콩�t�	�d	����f�%,���m��Y��n��A���t�E�ߥu>��-�K��Hw�a�)Q���*�/O�������o}�W���s�gқ,�u[B�M�l�0��d���t`�E�����ߣ��g��o_��Z{����~�Z5�l�0�%��S���oØ��$J#�=Օ��D�_/D�zD0�R�NS�#X�,��ƪm�^�?��(��0	�����gy-�����|oK�!J_ $gJ.,��~]F�0�Y�"�?����8�E����Q'COz}_���L��V���{����	5ͭ6�-*y�!��U�a�N�4�P���	׵��QZo�RM��*�d�� A�V$>�8-��//`�����2,�� Ѫ��Vn�D��cK����U�k�y��q�̝x�����)σIӡgʊ��	A����(z�F������^�������#=�}��j�H�L���P�0���=>>�t�Fӻ���#
��	&tD�|b.�2"
���6i�����pVV�q�X{Y�~�y W}�[*�[.��{���Y�f��F8�m�M �Qp$aKo�ݧ�����{�ݦ�h�\�#�_]����ʙ��Ͻ s;]v �<���.���3��r��|)@/r����`quG}X�{�_JЖy�8ED��P�kE�XGjk�L�i9��AN�ǿ{$:�U;ś�#�wDLQ;[��I����K4$D��^��r�u4ҽ)%��|�����g�OL��0Q�=�L0J���n �yh�Ѻ5�ɌH�C��dt�6�m8�Y�tTT&����BU��İw�&�^��9O�-X�UD��$�\��PK�N�f U�R�o��\e'㟻\��Z�{��E4�4R
`):4�!k�^}�[E=�S;�(��+���I���u�#�(�~�@��0��<���7nFA�&>.��#i�GAĵ���l��K�Ŗ�b���T���3�G=]W������X�ʉ$,��ړ?|N��}�m#��&��5۟�#�;�m (�7�US�<�M�4o0G�����t�B��rvWL ?Մb�Z�RH�s��x�w�z�x��MA���*m���|��]����G�A�/. af��ʇk��ͯ�z��E���a}5�^KԚv���{��~��ֈ���bp���G1[��܃�L��5�+ϼfJMe��d���T�er��3����u��5�m�雽�F�h0�b7�P��G$m�q�tfyI�����uP�\�=lr���tX��ɪ�H[�
�h(���r��b��#x}�(�8�6���}DG�G��N�`���"/��ֶ���!ZIx�߀�3m7�!�.�K�GW껊���q��z63�XW��ס/@A��A/ۭ�/sNn|�Td�l��[#<ެv��������,��a�7k5�Q�v��3|ū�ilp+�S������T��)�v|�2]��
-n��C�s��F��:�)�@yʊ����C�4$lF|��������iO>F����a�ے�����+8�3��� ?�s��&vm�X�S�W�c�ʇt���ϲgn�`��d�?,�o���ƾڟ��j3>K�%zs�`�{���ū������1o��s^�f��y�Q�7���rv �ܲ��G��`�":�Ĥ��[���-���u��������oɋO#D�@K��8��^��w��r8d��?)���y�^���ܱ�	��,��_	�ϗ��H�S|��H�k�j�B��K�v=�^�33��u���n~n��4�����s=/Rw�ɂ����}{�fvE���#Y�Fo*5Z��gr��n^a�y�����v��сQ3�m"�p�_���Rq�: Eym�\�p�J�qE��Nm����L�޸@.���N}s��roM&�;vk-.�B�D���gR��mi+����Q�6�ﰛ��1�y[���xg�AFF�TNs��!N�$"A)��&?��E"2����M{M��>?XC������M��Zq|���"�]�;ov��}_�o�	so�o��=��O��T��.uR<��p¥��:/�#��n�}aT^ضt�^�� ��R�k��๗Y%&x���m�#��ˣ��s{��ܑ�6u�q7oj�0�CD�L�|�umi�������2o|�^W(�>��+���X� �z����s]��cO�c�F����]S^�5����5"R�X�h����-_��A�jA�:��7x���q��ջ	eUr��0)�O�er7�AN�-WBOy�ވ+�"�ߥ��dK��� �6��=�y���a���}�qՊ�{��t���~��0Ӛ�t*��j�CQ߉8=�Ɉ��g��	TQ������o�-p���1$\b�߳��ș)���h���C��~�՚��;Y�T{	�o�,Y,�[=Ǜ��D������9� ��ǥT�l��œPoڮ75�i��T[Bz�	�����GQǱ�H ��:a�`�eȑm�e�qd
z&~�=_����Bx<^�27�m��>t�O�g���4%.�B�r��#��{o�.���{��#��Wkv�RȌ}�MHr��ۦ?_�cƳ�X`�I�����yB�����{��?�W��/�	���}��|w��g����v�L}�>"p���ǳ��qh{�g����»]`�G��Ae�:xW���iiA�E�)���{�L�k&���!|Ķ�)���,��*Ο�|�n�N.�@��+x�)� �&B���7v�1
ͼq�Q%&���[�� ��� y�g��|�<�򗀍��l>�Ҥߚ̻�q�]u76ߡ
]A�ӹ�?�	���$]�ۮ�fi����4�w�t���6<0�q0�
�B�����=��ٸ��U���d�egk���
w�7��+��ո��n�I����x��J��榞����i39�}�lk��ȶ�ĭx�(n�e89���»�ns�͹���#���K��� S���]�� Y�nf�8�f�c���W�[ e��;g�C7�����A3����;�/�Ã�4��������߿�~��;��2'��@��K���H�t4@w7�0h/G�yS�hZiZ�����I�K���n��=�7e����:��6�4;�́M���~P����"I������8S��EViu2�(��F����B@1j��j-.�� �M'Lo������%>f��1&�������}��1}�/�=d�|��o���C����� Hi�p5���j���ڥ<+q�;i�����?�U��[0��W7�Ov�9O��A;��jE��@c�<�Ҙ-y�>ֵ������wZ*'�ޑ/���}���[-XD��Jy�Q���x<3�
Y��`Ŵ������m��0�f!�]��	u�t�cYA'�M�C���Ϳ8c`�?�=�x��r�;��1���ZI��$�p���`�u�����ؠ���E�GV(�	�wu\�a�����#� \�Y8�al_:�����&�ݭ���}�}�Wۭ�f�i)�oaÞ@_�Vhn�;���b@�Ṅ�a�E�V��x��m>���H>�Pj"���D�so��Mp�)+��:IOdh��a���4��#c�pl�o֬�x�]T���$a�$.c2E_k��G������* }ѡc����A���������K�V���l°�f���Vg�q]Y�����琔���afu��`���O�%�5�ټR������8�����O[�ǥ�9������*$8b��2��I�b������3ݤ'S�^���u���U[�^y9ܤ�v�]L#%��"Ɠ�t�]ֱ{�$�C̽P5j�S�����r����_��,F	!~�&V�=���xj���c��c)�50� �ğ�C�F����f��L\jA���8e'@,���9He��S�`d��n8I���P|Xʔb8}��*p?���stX���J=�;�\1�]��L����h�A��j?�!�����ӭ��Y�m�fzU���3{�b�H������~K�fƑr��T��	0�,T���bH��C��K�� ,���A��ٝ���ŷ��e��p 87A�� ���TN�9Wyʿv�I�K�<zE�ȴ���X�:Ͱ�p�X�C��~�Ht����}�nv��a�SM�NPN4V��BG �J#=��T��$�0�箊Q&�vgĚ�}�G�����K&p�4�=��@!K0���C!�%휤��>!�ڒ����Ѿ�p�GT�,�ae6}޽ot�3O��Ŏ����M�lG8���4������3�yV� g�
�� �X���I��d�����Y+f�!Ì�|����ӡ?��j��U�(C���i�78�{���+���I�q��S���UAX!�G�P��6�\��_J�)��_���s)���y���x����u&�CV\̫��ɟ�L����1�#
��*V�o\���\7/�r읆!���Q3�-��q�����1�8$���y)�i1#��}n���Ni��<1��446�/���%E1��8��Zd>�H�qd�W��ǩ?5�8%rOv;�����}`��nʈ�Y[C'o��Z�E�
���li�x�,�d�C���i@����dO�HiV��J��Ï��zǾ�Y痥5�s��\]���H�'�>ƌaB��/M�q�����n� ��`�l���a�<��`������!<�	���i�������:x0w�D߽袁�O�Z�WpVE[�����^�3�X{Ɲl�z��R�^n��XV�s������a?�+��Muw�.��_�ˀ+��'3N�ɪ}��@�N|�/:���<�
7
꧶�OI�2�����7��h	�?d	_V��g�J��2H�>9\��^�&��\'���̬Fy��u�^�׼2��Mt���!7�0D�N�i�o�O�Ł��jIR(�@\u�	qg��kb<Ϫ��봎�7���m�XB�m|����Ƅ��s<0���� ���%��?8�������d���)��Q����s��aǵ���029��ӏ��NV���� �grjI=�˱ �ڦZ`A�Ǘ�8��zLM+b�w�4.kV�d�Ϥ�n��&VŢ��ghP��w��F`]�/j�v��o�V�I����Ao�/�|r�{@��B���a�g�`�~p&���Ԕ�'6Њ[SvƼH��P�b�|�*Nk"Jb��˕�i?�ɋ�����ذ7brK�j��Kׅ�=Z���K��̓Gw��'�W������jA��	��i�B�t�d֏b5�OMPk��]�BDp�69�*����V�U��q�Ŷ]�>�k��ėg�*�HΗ*\ W]6��|�/�'~Ђ7�9Zϕ9P�W�D�2O�5Xr%HgΒ��i����_�u5gά�f��i��*(��8���K�9� �X{]��!�ՠ�����[
�ʷy"٪>��TV������҆��lEw:��:����jr���tu'�:��qMa��=w��kg��k �t�X�p��GN�p�땷 ���a�9��M�;�w �׷#�vu&�K�
w�'ެg��e���1T�<��3��gt�4>�l.�Y_�7{�Ij,�P�@HE��NxOl̰'%��4|^�P���J	�B�f%��H̳B08��t��"ri��#{4�/�}�\d�(��d���{���j��O�8�,�i�n\ �������=���h��/�΋�P�m�p�6�&�R�O�x�Ja_�u|�ڠ:<���F�R�@�?^�ܭ`��n�]���
8�)>���`%t:~2۴��,z�lg��(̿�#Y�������b���v�.�w�����R�����Qߜ�R���t�(�@��I���]Dߺ���=О~��rG�8HU����e�i}��-�Q��8��P�%�5�(��� ��j��+�O�I<�,�,���50�z[�[x�$��z�JC�*�ɒ�mP�-A�+��d��{�3*dL�0�_v��-���z��T5�z�����uTq�.��K���}B{�O��.���G�r2�(MUz�������|0�G߬��QL�{W���&��ťBi�l�߹����Q���ҧ�M�7������=ت����tT��p��] �M���_i�����wH¹m�Y��%��"{�I����F��9��4E�>'C��BVC�T%���O6����]3���ﱷ{����y	��(cW�F�W��e�U{�'���G���}r�����;�[�/�o{wOýYC���Ga%;]G�M�C�Ǯ�?��)���� '�3�����F��{��!��Z^)6��=5-���:'�T::��D�.ɷ�3h�G� }�K[hݷK�#Ϳ_�V��A!��u����&]��R03�!?�:����%-'@�K�̾a�;��z�����F^\��&�Yj�_j��4���h]���Ә)�^����iYwvO�L�<n��~VV��ry�����^,E�!;��W����N�46��]��v��C��EO@�Ot�t����N�u��L�ب���ߓ��2�.�
���/��<�9��E;J�b����"�e����%�Vo��9S�n��#)�B�CG[�G�ד��]��n^]��7����<�h�/ҝ���&Ý
n�gS�p�x�߳췏'�ճ�=�q�aV�pEV���[��ǆUbt*ag��R���0������/+�J�h
:�6�s�<|�e�-�Z���Y��;&�;qL�����r�_<ω`�R�E�Zw���t����N�G��'�E�&��+�c��Bs��K�H��Z>
�`�o��=�Vi�٨>p��n*���_a���Ҷ��L��~������i�җ�n$e��J.����mk���W���ȴo����\��GA�oҧ�Կ��x��0
l7׃�������®�� \D��VX 
-�+��=H�8E�$D�?»��5�6��uq�Njk�
�W��S/(%A m��O�uJ%�±��:ծ_R!���@�#�><I$��5�8]��t�s���d�#�<�屮"��U��z�+������.p�^I�q}w��� p�cj�Jp^�K�P�D[���ă��J�V��-	ؐ9j�˲J�'�1������Mg7$�Reky/ZUj��Sx��D��Կ�)��f��0W����ʼ\��Ț9w&ѵ�
_�������6`	�����*�u丨	QX!�nɼ�,(�h�*B0�#�������z:�k �hȚt��\������m��xn'�j������ܒi�L��g���l�7���4gWO$��}�||p�;H?-��v��M��� ���_b*,o��?�v"��x{:���[5��V�;.'t4��,�)�*�������7yպY��}>tqS���H��ND�9�n���ۑ�UȽnyg7�ԁ蓴r{3�/�`o������T�W=��oůF�)��7i/D�8n�ڱ�����l�n���&���
���N;t|����+��T�Z�b#���G
m[���{c�_]'��\6�����6�V&	���ͧD�7O���Z�]�u�7Kd��Z%e�����}a�Ԗ�Qf��T������~���<���'�)?�^�b�͹/�!*Kf��w6���DAp�����zh�5Y���B�w�~K�Om���!���G�xh�8{@a6�$�T��Sl�&�Ў�'a��ထ��F�7}Fl�d+j�܆&�mZm<НC��E���Y	5��d/��������[A�f�x������i��>^����p�~"��\��N��������@զ��
��lD�*�.�	>|�7<L$=Nirii���m�� ����v������ͥ��o�)E��I8I'n��Hr�v&�:�ɒ#�+���#�w��6P��|bd��Jc6Q��}�ҿV@+�-�26���B�Wg]?�y�-7��\�	*���tqጹ9����Mi�{`�x"����d���$�-h��X�sw�
J��F���l�}q��Ѥ���ї����Ů�]�:G���M#S���yg��_&$�+QWZ��&νjZ��H�~N��5�HX�a��8_S8����X,��X�9��d˥�C��"w��\�Pw��3�́��lC�����@�!GW��m&绊�w W�Yw��[���Q��*;��(��p�$@���_�
Ӟ��59��GEᤴ�+��8�����%�����;]�����On�����c�Ϟ��/�]��|t�_K7M�?Y��g�9�/홭�`�;�W�W�P��yԚ؇�7%\�w�'��}�4��x�����Ԓz%M~�AP9��0tnP%ȡ��j=�4�i����)��x 2��h���P����N7HJ0=�N�ZoÍ����tnsq )�"2eH:��
�x�Yp	�0�����o�t�VRdh��;V3r��ry�􃿶�E�]���΀sR]�&�K�#B�d�j2������?�`�z �aX0��3<\͓��`Nʥɵ!]<W��;�|OPL4� ����s�W�B���~2j|rvX�K*��Rk����.c/�3NQ&)y�.���R�	{7G��e���+��"��%��=lPJ~/�@�->�O�W:o�ˠ��z_G3�'7p?����ó�,��ܚ����3��IRh�F�Ћ=p�"��m����[x�"h7�50&OEL�#A{��0���r9���Ѧ���W�� ����$K�F^���ܣ�(�hĮ@fiY���8M����r���=`6��#O��Yd�5�#tܝ3tQٵ Q����'�@䳇���������`���L��0�wN�I��jk���2fVA�,V=��}?�N���A�;�K����`T���=YYB�шro/0e���0%�8�7f"�^2��u��h�qS~�ji�]����w͂���/α茶Z��| ~�����Q�:V+��g,N�.Va���R�pǿ(.�x�2��G+��Q�zi�e�n�NO��'T�=�&7�{�!�nL(��f�I���%�Lo-��\Ҍ�6گ�t��W�ָ8��R�8=���f\���Q�1���h�-��-(H;\�G�:]���ٱ���;�#Q1OK���M,e]X"(|��=Ĥ���,�����1�_Y�I\��������R\�tl�f�t�r��G�����Q���$u1�l ��y4"�q/�M�"�h��>K����~�Y��/�n�(d}�iΰ�bbL
S/R��l�.R��Q����N�l��(5��F��wßcS4�5��/���_R���9��,�R|A�|LK�Ǉ�f��g�����=�'n�I'*�M����.]L��Vȩ��$;����
{X
"��*����VǪO�>�I��U�)L�����d����|���g��G_t�?O`�i�����vPO/�c�]�9peO��8��?7�����!X6m@��]"k�<?�c��qˢ����H<�s	C���w�YeW+5?{��D;����2����4�XI2Q�oL�'Ih��
F�m���l���_����3Pe���b��*I����E��yaF5Q	4��O`P����7lu!fݦb# ���%�ɑJ��
���z�����QE� �I]&T�r��I
w��m׎\y�q�w��;]Ƕ�^��<:A9����ܤ&�&4���{]ဖ���jǷ�Ԕ��O�S�aK�����Օcb�{}U֋���0�N���p ���03O��֊"�,�:Z�K���tӁ,�CCϴ��4w��z�/��l�Y�@w쮝�z�(0U� ���h��`o�Hر���V�뽷���Gd��x��I��^�H�ڦ$��|?�{+9V���m�Дh����e�s��Oe�r�]�I�7%.��<44�B�Г؉��Uٕ�.Q�����ͱ�HnD�Fy�����x4���Ҍ
�2!���ҥ4��֭�ї�H�R�����m�7��{��X5,�O�#s��n� z��2>+��i�80�	��ֽ�Mu\	�mW��^n젢DG��~Iq� )�q�VY:����9��rOb�j��}G�ǐ��_hᕸ��L��sC�wy���RW����B
���XKvh�+�"q�#_��C��梟�TUX�#9��Yr�s�?5D@�:�^iV�E��qh~ŧ�nت#SǃV+�)ޫ&(A�R�<0�2*wu,������I�4���T��^��t*��ȸ�3�I��Z�H$\�Pf�?��X��\�,P��ց�y1��;�Q���K����.;�F�;#�*V�@_�p�H'h2�%���T��,�l���x6��2�]N����m"cD�/����>�낌j~�6�Q�Lw������h���T%�q�h�u�	1т�
���.$���ˀ�fp�ki��NѝP,����1�Ϋw��uON�S��wت|'^M$����i���DӸ�E<�K�1���������*MN.=�_��d�A.��I������ϥ���{՟��;��J�\z�� ����B�|��~/�gG	�G�}0�ǖ�����sLW�� �{��5��GRDO7�9V��l9z�> ��6�~uw����l��������ZXa�h�ޤ�`ٰU�o���D��������݊.fR�;�[X#\�lZ?������^P��U�K���kq2]���������r���Qұ�K�^���OD}����X3��L8|���ΰ8�m�;�5x����ogN�]��H�$T�M�y��E��O}�A:�"?���|x�ǖ�P�G1�~8�[, V�쑰9<�F6�؎�O�ϯ]WW�B
�!�\?�t�nĹ_=^�}4�^c��G����ۇ�����_�6��s?��wv_�m�B�	(��~ڭ(D_�����Y�}U;�.���胦cn �s�a�Օ��p�V���Z>�,�^2E z����N<j:�����P��o��'⻺�q��`�8�T=�-�;.?�V��$Vs��ҼG*}���И��N�Q�Y��e�\�49�������x�;�[����{�\y|֢�j�M�������U'�V�F�a�Nl)]�_��H*�^+T�%�]�=(�s��d}��o�s�SW���f"��(��Tz��+ ���O��J�>咀��Πp�M^:�T?Aju�rǽZ��bݻ��c��]�ԈGQ|�<P�����cݠ0c���bZW}��j�7���=��Yt¬�Q���֍����3�v8��ۗ��G��w-l�������eqxM$N�p���� ⽼G\؞�l�u F��ri�K-���O��5��-h~6��
�Zx�eJ���*������y�w�'0V��◗����"P�t�Z��<�\��u%�D���Bp��NoM���q� ����k0�c���
F�T�s���/�[���Z.���1�k�M'�a9���>�[�S��륣/�V�y�U� �s��7�x�/a(��#�}�e\�kdJe��;lm��8��.�q��fu�5�H�Sf�,r�;13IJ9d�/�j4x�9)F�k���tMKܦ��s�X&���7��ɯ��)�pS_�F���Mz(��0���/�5ݟ�A�Y`��"�[s��m��Bw}��$�A�S�ޏ�%��3#oi{[*\�}�,��:��|=�;�����~$�+=�pڠ��������~[���˥��D`�� 8��{��V>5'Z�y�76���%E����8�$����
�'\*���f���3F�ӹ)�#x��ceq�y�]>�7Sj����Vzy���=�A���yZ��"3����LER�����'�9vh�Tg�s�|U_�������[<��#ȑc�6��U���r�<�n	�"�B���6�
�ç�����|T����wHH*%��C���$��1M4�pO���p}S�~͆r�ŷ��;t���
	��;��<Q��
̙��'���FzV�/u*������q�/�մ~X�(��^Q͡��^H�`�hMzu�3L->�/���KD�����v5��-��
��^�DOelԢ��+U�~y��s�0���n�� A>�j����|4�<���X0�vG`z ṲJ�`��Ð��Jb/�g�@��ͻ�ߓ��f�4�9��������+3&I<���^�){G%�0P��vEٍ��ۀ�o��:�0���K�i)��F��
��U�LI���ՅNL�,㰙�J�cSȮUe<�a��8&�5~�I�9�y���{̑_?�Ъc�V����k�قi���<����
�GH���z���s�H�®��؍[|�┧}�>,��r��P�hFђJ�'t_z}����	9OӉzrA����K��1E�g�I�
J:��'��R ��z����~p��%��C)�-ӻ}��߹��?t-��ތ��)q�H���>ȭC����4�R��1s�c�r��B�6\��{���@$ɣ�����.@z:����)f�o��g�W��43���Z����YJ�oG�ئ"v|�?}�th9��h��/��OV����z_���O�E}o�J�t۬���������[A /�>��p���sU�{A�r��`�h��$ۮNj��I��ZEwr�&��vwk`F��[4�-l��s�J�����s���y�N��	v������I_C��xV�ՙ�0�D�����O�ER7k$y�V���3��
�y�Ϝ��՞
6F����^�z�wF�5��ⓘ	T�y�}��7�m^M
��ʩ�۵��`�p!$�<(9�;;��A�$�l��'��'�ߘb��+})���º�����`9�<5�6�����8;N�gP娻�V��E��vmܘ06�A�H�i�#F�C4s����Ōe��ƨ�zG�h&'XN���*�9�a9�.X7z
�;BD^���_�/y�8-܈v0lC�"G�g��,0
7����SM�k�\���V����V�������������B�rq`�妱��I���(n��p'��u�����!T�O�8@��L�D�p��k�J(�]&�/�|����C���I��'��a����nF,*��/�n�x��;w��ђ����8��j���e��<��OJ��}�ٶ.���ʨxY�����M6�^ ńtX���|������, O�/��bLz](�VԓĨn���eON�:�R^]�h=<�e�[���R��t���M�W-xE\��]�a���`�Xːn��&��L
���_UC͏��j�������oQ}o�(Hw�t
H7Cw	����tw# %" 9�HIw��CHHHC�H3�٣�����7�k��a�g=y�k=k�p����`�X��V�b�}⧭� �P������lƷ��I:#*�SZD���Z��)Z�`���.��b8����k���A�͑����ѷ_�op�ō��ln�u�"��0�\*��9��Λ�>�m6c�ë �'���o�Fƨ��=i�wÎ��]�|�s<�4��Q��\�O1E�i*�����`Z7���CA���f-����D{�L���ĥ�)���~ێ��-ߚ�WП������<f��onO�L�OZ����"ʜ��d�گ뭂��'Q�n�B;�*���!��A�'m㺔*�z-]���
�)��tx�u��8��1����m1B��b���#�>׉�����Z�p�=%f�P[��"��YH��fh�^l���+Yx��92���e��U:9^�q)ِo�NJ������I��Քh�Y	�0_�?ɉ�f����a+��˔���b�z+o2-CG���+���&l8.�`�'*�E���x9W�yA���j�7^ES��F]	�K�cu*L^0�A��¨�B2�Ϥue��{�VB%Tb:=l�p=do��j_���]wv��j�H^��G�`����P�qx�<��˦܏S�2�ђ���O酨��[�!5\������U��<�7�F�*�R��N��M�3f����5��P4v������7�����DiL�8�O�W"^�v�7�䆋�� ������Uo��|#�~>�G�FnL�����A�f���������@
���S�-U�X��ͷ�w�G�Fn�w
�Q!$s���.������ɼ�5L��d��l�+��G����P�얫@�-�ܰt��!c�J�����"���1C3��՘<Ön����K~���L:@-�s�6�Ow6�f�o��F�yv�I�� �C�׀<[�!>p֭�����\y|r>��jt��r�K5��:/G�+F�B���}�W�PO�-�ũwSE�cl�`��΋���GVA�3��W�S�Z���@���5�ikl �W�Q����nV��쿖p�x����j�����ͤ�{� ��q�꿨�l��,����U�i��5q2Y����E���%��+{��j�M�#�pJ׸C������,K�'
��~�)�>O��"v�ڕ��%��1$^LV��lى<�X��.�:��>��iu3vc�g�W6ȭE;�D3�i��VE���>�7���K/�	ӻ;�3�/ԏ���X=u�¬�ꃟ(���Q\��d��q��z�U�-<�J�P�->�tOK���5e�D��\�!�� ^�$���*��3�kUc�]�3�S����͢��r���-VV_�_f�Z�d6k��@�q[K������SkH��?О�'���D�3�{��������M��&#2F��"2�_��֋��i1��_�
H���r���H-�qj{|���ԴEA�1o�F��Ǐi�Tz$��`^��K�x>����8J�~Ɠe<���`���m�LC�;�@�_U�l����Xo��>��ۂ$�4��}��-V`s��v{w�ߑ̄�j-� ��jHz�k��q�.�HC� chd�w0�R�~���o7�Z��96�i�i9u��V�N�C��8�N��v������&��|��;���R5�[�^���á�����q��U�q/Z�$�><m}���� 2[��_8���i��3�?�Au���� ����I����jB�z,[rg������Ϡvv��rJ��jS�qۿ	��`�@���f��cXx���g1��Ѱ����;���T�Е$^��d�,_�K��}�s�b[Cq�G�t�.�f�wt��tF`�`�Z�� �����N/]D�.�U/�=D�(_��1����(���8Y�;���g�{L
��>1�?�6�Q�1֘��AM6�D�v��e4,��7�, ug�g��~�E�ZT�p �%n!��j��|_M̮=����D������9���`�翂lI��{�L�"gɒ��4O�cOd/�Z�l���_8VfV^ַ�od^�ōq��#��f̈́4ʔ���lMX?sߞ��%�yӿ0�؏��9��(T����H���c�� _,U ���K[�ߛ`�783p؉�J!!{-,eo��G�g�J��]���3no�B�Gݭ4)b�0�Y�6T��^5���P����)�y�4)<yO���q���C�m��b:�NO�;����g���  1�$F6�?�zRz N�z�!ہZ� �����|*V(�������� �"�3B��n���o�`(��9��U�y���@���U�ZDz�d��Z&�n7U��������eK��B�wP�'>�{�k.���E�.�>.���/�s��pk����+P Nt�K�f��YFr���q�%��[��<��@e�E�X-��?�s4���	������-~�>��ү�'y/?��1��3�� �N A���ɂ w[��>�C�Mƈ��u�����Hw~uz��L�J^~R�X'V�d����K����-�8��Eѕl1/�A�b��#ݪ��N"�҇B[TO~nR�1���CJ�~6�����8G�ϛ|r����.���b�����'/����["��{M2Q���#J�p�U��2,x!��h���Sř>?4�eH��z���|����6 �*���)����:�m��Z�Ь�������D�N ^	Y�%~�*��k����8'�g�d�J��O�XSKRv$*Lmo�Yt�ʟ�|X���"�v���eT8�����I��&|(�l	T�A���t�r�x�-�=����ώ��)3;�w����8��ǥU�I���-��
�I��8Ǆ'S~���3�<���N�������Gc���ƧR�,���B����wL��dYg���xy��jI���U'?T���.�Z�o���s,��f^c��،r���˚���ȕ�nI�;/�R28����Z�1��W���^.�d��M�mrp>~8F!왕������d�n;�D'�p��iZ��������t[���\�\?L��	����r~��V����x�������������ר�X���}ɩ�F־�	
!�B�lR����Zp��`[��` �Dϕ���ۯ�y=j"�b�q':��7,[��Vab����1l�^��@�j�{6�[�s%վ��p��H�⑱�����=h��"q��@_�s�0'�	kw��O��j�0���A+h�5��3���>�i��C�T�Ot��k6�Ζ��f��Ȉ5��Ơ���ZyA�ޚ�aY�e�a'D�r�")>���$�ZY
/]�o��Y�Fpm�����1����O4Op�=O2##�*�_uh=p����'�g�;���L�\�N�)t�u�c�+Ӛ�8�+��ఊ�]�h+�����9d	i�� g���( @1�Q����Eט e�I��Phoҭ$����[u��>��Mˇ\>�3&s�s�U�+Bsu���������9�Hax����*`�3�aD��Ŏ
7t/!��k���8z��v2��h��l���mڑ�]zV7�������9P�7�9w��kƛO�6�,����OI�e{��&r��[��a'�']�وIѸf��5A2�n����!��߽5��F��&�k���&�0�l��>$���J��|�_��X��S2iȋ��yy��Ͱ��Z���K�U3�<�/��:�,����y/WM�B�I(�#OvX�}� 㹗��t���/H���S��z�@p�;��I��i�G7���q�}�#�L�3��v��C�7��wo"l����Ϸ�7�<{[S*[��ᜋ�(u��	c���ol͉Y��" �/��, �j3%3�>���W�P{}�0"�����7IY\����#a�= 3�M*��o>!oc�]�)�Z�{��U]��a%�x�$F]����O��9�6Q<@��0b>��'�gu����T0!�@9cJ/#Ղ"���1H#ǐ�ծ\n����T"��s �����!�����=u��I�N ����o���a��l�Ʌ���u������O�oiu�8H���Q˩��Ny�򀝫�U�	��
�g�Q퀱�P.�R��hS�GW�gDB�h,_]T�½Y(i��{@F��8��t�46�t�꬧Ȍ܃������t��7�	d^��-���eW��x1��/۵����F.�����6��0T�,LL_:�|\�U=
��_�v՘X=�s8j�w�!��'�*��*�t���e(�X������r���x�̚4Б�	Q�������!~a(+{��\Ư<�4�Q���`��"�[?�/n�%�l���O!s{z�B�у���NMO�%!�X?;��Kl�B5�h�����{&�F+r�wIk�����&`wL#���$�Իh�`N���@%�&��?"�!d6�����Ї��D��6W��3P�`j���0q�c9����h��ZRr�=Qnu^L���S�t|1T�].4z������}�q��|�#�\�������vC��~K��"V,�0k�ver|?lŝش[C��ߖ�g:<���z��ë�i7 �=_�ɴ���f��,��	�v�<6IX���ʕ
�i�Wv�ok��p�n�.cnmr�9���1��A҉��]k�=H��3��jԷ�EE���o9yb���Y�5$@\�� ��򌦋J��vL;+�S�ʪ��kk}���fJ}�)�,���_i��P��#���<.��W,�N��ޖ�Ϯ�<��?:�pH�Ai la�,�0;�nR��9����X�����BUˀ��e�?���ι��D�K��bA�����	y�B�Y�`�S&�_�j+~,�rB�*cB�b)�,��	>��<�t�R��~���PP.\^FVY%�@��/���1!E<ĤI�� �2H���rmږ,�~fn��]�+b7��4>GX���}�i�������3fn�R����Y���ف�������%IP>����w��f�Fܟj�q�`w5:�&{�%�^h�r,g�T�tr�>��"V4,�~I��������
��<*a�r�m���P9��:��q��	�|�@�t�?�[\ZY�E�?�̨������;�t�ďhVP��w%�S�����//$vE��ʲ��8	X"9	&�@�&� !��1�d�zt?>��>���@n�@N��{��
I���+į���XM]_�y��?�Qy���j���1��T0��r(E��������p��y*�@��	�Zf��_'���>���ST�Q|Ī�����`�ک�)gC]���<���E��Ma)
�|@W����i�`��]�o�HQK���_���՞|z��R)Ëw���'}��MBx�ђ��Hn�4�q�B�~���ƍL6�y����d�����1��U{	A��EC~廩a\F�Bg&KƥCD���e0�����ρ���)�b&i]٨�� `��x�î���rR�בq��is�������'�d8�e[� Uzw'���L��e8n�V�/��Pۛ�|�?��}7�!#BB�!f$���Y��6U�?��ɜ��ګ�áKp����1��;pf��.�4�f߬�&�,.�I�4}B=����w�0��I̞�Ri�>K�V�'1�z-���$�l;��U�;]���"wt�;=�P�+ra��j-��'OV	�
9�H�9�}'^ �Թz� �ͼ�D>q����	���!w7S�����v�д"@��)S�HF��w{kj�G`6Mt� �Gyh�9S{�]!rD5�8�`UR�SeU��v-	)��Ҁ����h��u[�7�Ӡ���J;�p�g�H�!�g�*��߿K��d9�_E� ��G�Br�����bS��dk��"���ؙ������Ã����c��ޚT����9\�����Z�n�W��KHJ�5ic�kO)��O����� iH&N⭽����I�}���iD�K�e�=&/��A������x�~=d��P���L�ga&���~j�^N�d%��0,��@1`�
��<�)���4��������'eUNS���F��m$�U��U��2
 Fy�L�>/�l��CN� O���P�G�]�Ve�&���dI��M�%���Q=��W	*���
������.�x�|��^�1
�q|��Cl٩�TN�R׃7�����Q�'p~Pv�T��U��7� `�g�=8"F��|�;s���ف���Κ5u��γ�s>j�aN���{?�ݙCܻ?�N��*��X�@cy�L�=��,���<�����ء�03��W��������I�N3
�!��D�JNg�~׬��c�j��(���Q�(�?;~�ܶ�B��s|(�����eh*�ͭ����sb�ߓ��r���a(��7X�&����l���ĩ�5�gR�U3�>w�'/�FW��eV�2!�;��H����u��?T&<P
8�χ&��Me�|
���1��k�<7>@J�|����M���KSN��R=*C�}��"40$��z5ED���	�����6䍢_3K�-Kgs�.^�X�c�N&
�rMk��LS���V��c,8<�sl �Y|5\��������g���C�t+7��k�)
J��&ذ�[�"���LOM���x!�Xċ���?Lk�p6�.��)��@��� �a���������*	 gȓzm��^�߮k�W{�0�B��wʴF��N9ryW�O�,�V���a�;�9z����Gf�Q"�g�:��˻n�
GRh���L�,c��Zb�oB]^��u�F��x��c��.����Y7�U�{�ߦ���?���/���Ḳ
����/9�{�!�f�Vq���I�K_9�]��%��08�y{�-;�����PD'-��K������/�QĀ���6a]2�ʣ�r/J���˭ّ��(|��7O�������=o���Q$�_�(�*���F�ڬ�C���{��wv�	)�?�A~�WSA��O��4]S��j�IB�{XD�������	j�_w�o��K�YV�~�lfqǇ&��O�XX�B��	A\ȧF]��.o�8����*h+��s}�=�0�/�t�3��_4�(V1Z@�ūQr�8Z���(�9e;{��K=]�?�g�����L		�r)m��%3�괌��6���O7�
S���rîb��р$F�ځZLP���K�ꋜ����������� �B�
�p�M�h�����5��P=�~�W��	���X��h�����>M��� �1��w���I��x������#�'_�����j-ZC)BG��b� &�l�Ɋ�p�Ƴ��+[���S��4z��scSRTGGw���+���Sv���L��`��IoK����;b�u�L���	Tg��b�wS׉1�m��RB?%�@ߚ�����ob���ۦ�\r�����<>jꦹ�!L=�7{&�ge��F80���2�	�����_Gax�J&N������ �2��U�Z���D��z-/Od�pB���,��B�ĕ�Kbm���x�y�Z���a4���UVh��P2�[��%dR�|����֫�r>�a'�>g�);�;��"U�:e5wN �Sv衣�9���И���a�6�h
�ҲN��a�؄R��X��6��d;6��j�IJPB4$3F�7c�g�&�����B�H=���n�PZ(���C��]�wچ���{�(g��5]��/���������c�#H��P��B�}�l��ӿo�լ�)�:h��M��ϐm_��P�c>r�x�_��$�>[̻����d����%�X5i��(ې$4����2Rw����@p��K���|��v�v���}^Ӷ!pE47?��b�(!2��$�w���8�-y	E���k[܌?�F�̏������ /d+����E׎#��(�YF�Q�;bGz�4/m�R�w�W-Ԧ��M2�it"�{�#�,u�)qS6qS��}��n���h1��/��؀�����ĔQvt9�Y��MN��'/��W��=@�X�o���k_jN�E �s5W���e��9$�9�W@G�"���h^�c��w[��C(B�i�uk�I+�j_�vl�s�W��Z�����:E2S��u$��?�$����.B?Ҋ�IXlk7��w@Dڧ�cL�Q��(#���@O�����������f�N앎R��XEa��z-���4�j��������_"�̸B6}r8�1us	怹�]�Ltnv�����\�b[>=cG��@��cщkx�dSW�(2�s�<�:�A�$?%!�C�Bip%\�]H���2��/��������o%����D{[�42�i��#��K����ea�]���b6+?rO�Q�ƨ���'�{߷��_�-�d�A.�r���V�rI��ؤ\V?�M��+����H��Vr��0��!E���k��Ko�s��7w7�
�U�6���5U`�KU��^�{ܣ��iH?x��)a�\s� y� ㊒x1[�u���g�	��S�iH Uv{�_�Z��=���v:�3���D�
��V�p%*���%E�M'����^�ױ��M�v�C�
��+s�}��f0K���^ϣ$!	%q�<���B�P��	Q�F�߿e�����_6&�� �edυ?�cM}�"���=�O����`��06�J~�����\�8�,�48Ϳ�+���B}��}����ؒ�@=M'�$Һ��	�dpb`�&])�c�h%�[1�Ѣ�c�v�r�8�&���`��}��ḅ���	�-xM{4��KLɘ%WW��g��-�{�l�r�04[��K���d�o��;��8�\�!79�Gq���#������wR3�5��kpb�颖.�s8�~G7��k<�g��M�:��n����_��r		=��p�-楪�*f�ZDF�
�͟�C��s�ϬZ�X;�fVƍ��� ��7�E�/PK0�_[15�zs3XN��O�%��Y��=��S��w6e�"�DI������4%-��%�h�]�40��ԓ��H��4��۾@P�xD�\�F2ED�`%Ba�A���-��i��h%MJ
@�$�-�5�ċ�L	�u�ʨ�/�E�Bt��l�$^�^�����w�����ݣk�Xv�j�M?���_�dM��P#�Y)���?Ӵ^��J�;b�)��\��&f�1�:I���t6����:���	%Z��W3S֢M�rg}����]4)%�H�b�t�����東.		(�&���>�i��rx�������U����5j����؁��JQm3�
��
�=D�����`�q6_��'�P�+�o�:�Y���Sv�9��E�˟��s��k��ՍΥU�L�Ϟֹ;*���f&�vgs�L��~�5Nb�p3E��\.�a�u�����:*S넯f3���kԍ9�]���Ab����;m�X�4;pB��M��,K�lf��%����Y=h���n��U* ���R���_�[���* ՠ���h/;��y�C��[��^�AJ��Դ�T�\p1C�i)���d�Z@����_�r�M���>���i\�H����fm����u�+R�����m�=X=j�i���|��[�!Y#���76 W��?�����<���w7�3M�AFm�C�Q�j�-f�A�-�u�/����릫c��_$��+z��G��NkX�bƏ?5��$+���0Xj�wz��I�di�����_�߈����l��h0o��z��
���d���w�EHے'� �2@�^g��T�>��@���3W��,��.�6�ݶ�:�,rY�"-+@/\y"$��ȐZ��\;��_�\)����>���� �Md���{8���n�2����_�	m�w��-�M�VED�����cA�<ܑi�=����#N^i�?� �ě]U>�L�Q��h/��`���Mk���p|Ih��'c��a��n�锡�,�&y�Q�J>�0����:P�en⸇�wCes��Ƭe(�z�z'A#D:����x2I~��$�n�`����D�<�;��w� ���&��M�og�J(_-���U�$�`�'ȁ<ҋ���ߞ1N����y���g��2������3�����-#���?8�<��ѿ��Z�>o���c����j']�{7 �1�~�����{*cZ�{47����H���`5^G��,�&����}%fNO����0�4�f8p��s	'�C�;[�ӟSAw�m~S��J���_�[Ƀ����ī݆>�3Dt��^T��w8�{��y�݄�Rk�:�E�_�C6�|H�n�(S'V��ܖJۉ��������F׋�?�_�L;Kk���_/ ������©��f�2�3Иc޻zd�S�[��9G k��[�>aer�k�w#L�E���˕|2e?�ta3
>����g�A��4HQc�N"��
O����[ƴS���v{���'_5���wϘ�~��l������R1 ,�
Q���2�'�Q"���B�_�?2l%�����3=0�)bQ3����h�Zk>'��5w)Z��㊮��VI[�QK'��ZXulђ��8&��VUp����x�m�`�
.�z��پ#������R\ʻl���b'�s����gs=�ް�׸Q~C��ɦ��C+,ˮ���(<���������eD���4��;CJ4�O�,��K��Ǫ�ΫFƛ��#!�g�%06���i�^�н�3���y8����l�T�堼�QU���SJr��ZB�YBJ����pʧ��\>��i���;�h��+�ܶ��2�(wDNm�y�z|�Q䗈�&.�Qv�d0�1���h`�Y������@Q0'�w��zv��n�� �s2"B����A���7UBR�g<�������ʣiY��Vr8#ch3n��tv��>�=�&K{$���/]����]��P"�tR��W��;oO
���7_k���1R ���m�<�����4I�zNY�r�l�rxi�xf��G�/e��O͡�q�fj9��0�R֕�ܶj���[���MX�v�	)��8��f��͆�
�^!���S��w'�ċ|�,l���?k�n�vkxp���㐘���'$�g!B��)�������m�m�;����^�:��{U�qp�MKYp�y2(vh��*i#s�bʡEJ�a�/�}��FLB����52����lR�'��ʐ�O��>|^I��뭭$џ[�^A���6%��r����C�,�9c�(�ׅeu���J�}]B0���X���nf�aA6�'�j�F���V����9��a,��JK��Q����7+�����΃1u��d����dt�2]�M:��_t��zHfֲo��r@'4�����b`�((s3�\��>����yI)���>�Ө#�c�~�_�����������@yRڙn�u(!EaŚF�ed�Ĵ� ٢ ��n�*�k��pƤ�õ�-�����j������n����ŜF��J�q���2��ؠ�Z�b[���y)k-�ma����#	mW��6�=�!�5R�
8�3s#��:1�����O�XK‰��XY��fs�bpl�x�d?���r_��hu���䭚@�Շˢ��r#c�}�v@��E}8]�o���(��e|
G8��V���x�:{Z�^w�]��w�(ReՆ�6���bTx��V����k��Ŕl�!ߩ%ܻ����}5�#��3��F�ɡ��N-8�En-d���K<�z �ٷ���6$�t}�Of�M�>|Ȗ�1�Q"��qF��Ʃ���ȁ�;[u
.�3��aZ��c�u�}��,\�ջ�WB��Qjj����
~&�B`u�.o}n�#݊�պ�4{-���U�o&)P(�Y�-� <'(L}kv1��0�c?���� �O �4�~�e۞Ĳ\��o%����Y'ݷ�v�AJ��U��?U2?�j���J���P��X��-�.���� 6t�X��ڝɬ��m�:�wZ�
q6	�U��"�/���\�2^b���F	
�2�;�)1��:���H�?QP���)@�I��j��q]TWp�+%΀�=f[O8��m���Q�ΰ�	�w#C+��&�.&cN���N�+�_�d~�~lf��ЊH���{Da�W�8/*��'�C�\��=EK?�7���*�r�ў]�Dř�@6w��	�l���4s�{/2�o�e��p��8E�:��c30�T7�#Ye%B*�9��2�o��U
Ĭ�{�e4�#�����P?ӵ0�/��� ����Y�Q4�c��������l.:<����<�� �j>;\G,^a�9�T����zyκ�N20��V�[J�*=l�#�V�J��U(�P<:4,��c�2d�gO�����\c�r�����i#�#�&�$Q��x���oƁƓI`�� ]�՛K3 B�	��U��ӗ�vN��g��׏�5�����I�d^�8���NNP+M�K�P>���Bd�3�ڈ"ϹKzz�w�=����t�^q��y��d�</;��c���/N����/-cW�-�}3�"9����=����Z�=���/�L�K�����Q�&i�r���ڥ�����ROw�
�S �@���W�b��(�f8��P:��lV�CRB�!Fy��z�U��r��:��J�W[��dd}�������$gӟol�>�Q��&��΃���hն�e�w�!ޡl�×�i����Ae7]'u�H�;��Jz0����z�Z����ƙ�2 ��zD̑���Zp�H�B�,b_�+�M[xc��ʪ?aj<���bvO/G��^9[�,�j�<�Wi�т����P1<�n��!(�_ܩ��qY�����.#��쵚�G���n2U@]@��(�dq;��Ul0P ��(�I�0��xH�@�*�����Y��{�5a�]M�2��^�^� �l�R%ؓbK��j]���Ox||ak����u���oH>IGî�ĝ�ƛ�I�]��wL��ϻp��M�߄b3r#���oB�B}����.c">�"R@E�F�P�dݚ�y�[8�����7�v���E���QL�UZ���w��܄��Rw�������OU��Sg�{���.}���J��d�?&�Wh+�kEA�ݢ-�M��u�E��������nWJoڪ�x�$�/��%��Z#�~p�����\
S�G	�sU��Z?�/z;5>�/�̮"�ѹ��-�qdu���X�&YI�,qz����"nz5�BN�~C|�Cń��ǟ��{9�.`��)
�q�Aȃ���܂��h���j�k��Cò=3�Y�߲��ݪ�j��c��I�7�d*�/�獲�"�9��H�%��Eђn��3r�W�4�<W�|�"1棖W�b%�Q��(����M4���XVW�b6�X.f�x�g�D��w����&FF}�F�HU&%p�q���\H������l�s;����k��5�w�_z����e��Ε5t�?IB�>��2ؿ�	
�H�R<�Nبe�q$!I�2&z������P��^�P��Ic��Z�7���2��i�fL~�b���a�� �M��Vx�@�|E��h~�Nz��^]�16x��g��jb
	Փ���Ε����kXs���4����0�sޙF��󬈕�����Z�*Os��j��]���%mƆ���WCPq�a�T�R����J�����\�s*��r0��w<~�o�����j��E�f��_]��|�����C2��s�8XX@�i_�Bw���Y��#�2V���]^�5`��龰�4
B떥o��%�Y��Э��Qux��p�Љ�5���RZ�Y�˻L�B�n4p1�P� �qQ�p/Tc�x��u�ty�r��^��mؼ�]Uz��|�����
ǹhM���9�����-q�t��)+�;ƨ�3����)K�jN=%f���wj���	�<�s�I74�r�⒫cj?`����$�o�Vº�L��e������{U$>H���?�7	dy�j��X�^R'��T~���FR{O��H��%�WΚS��y���~8J�������k���E�+XKN,���p�ú��#cY���N���*��Q��ڔG�f��Բ�>��j�/}EZ��T�$w��O�/�mu�"�1<�;�v���L]FF;x~��eg E����,�;��K�,��ʭ��iP��F07�IRO��$6X��+��z�E�hq)�i']�Gw-Xn?�|����ڇ�����ۃ/�VE��^�>�x���IN+��X�2�1�����HJ?ދ��Bs߼�VWJx���U��̷�d����uX���VP�1o��r�ŏƉS{	�����>kk��b|Ool
�EL�
9�'�V��F��:��?#qX\S�ξ�,�B}��w�"���O�v���i9�W
�A��`(�]��>�t4W?a��cB7t^��ôv�/i���C�7�-�3�|@�����>��ٵ:}���(gQ^�2K�m~���G|궖���S>Iܰ(���c 7�< F�e�@@3m^����,���p�_b(�j;�:�%�N���^=�����^���_SX�I�S��u������-�<k�11wY\-���dҨ��0?����ś�	F�Ռ�A���ىgL�M��I�3'm�r���y��>��}��[8�����ׯ�CI�ث�S�)Qa�����/����}���H�4ÚF@"�&�y�gd��k����g\Z�h��$_���7m�Z{G]_��7|���g�w��5t7~p�Zρou�%��i��<��`��o����^;8n2n��K�_����Ƀj�Уr#�]��q��v:<i���7���ߐJ���������f�M�á���A����U��ˎϟ�<n̓���-��Y����Bq�;��P$S�g�g4 ���=�G{.t��e�֙�W���W��+3bJ@���af��^�̓&=���@ǽ�}�w����5I�:x�ks���`̔Ѻ��2�a���S����94G��+�]}�ƛ�<����A��s�T]�p2i���`��3��;5،����VJ��c �V�=Y����'��:pJ�o�pq�}�D��&2V�~�����?�`j<�����M�N��]o������s�� �Ն��؁�k ���xd-�A�#�;�e��o6~o� �k>�1t�C��^M�M��$�ϳ�+�ަ7�'�L���U}l�q�zO���u,�	y�O�;0�p�ռX�i�?�{��eM��ҍK�D�w"hJA��ʾa�)����Rt�jC��s�k�j۞�mm�սQ�R4��.2Om��x��yc�ϻ9q�K��`<�	/+��67Bb�Ĳ�Л�c����A��ur���3�f�QI��B�E}����=�fA,֭g�W0j������j$Bl}�5�s���-K��[`<Ў?���.�5�q
ǱB6}̯���sq�H�%"���q���`&1L&/~��A;�`�b^��e�\\9�`��������<X���җ��<�H��'4��q�&���ʹ4�^{�e�1o�ߣ(=�y��� ��å,�JJ���J(��M_pN��Ϲ����p����m��:��4�]�5�����S�z�`ϣeQ�Bf�+W�4�̜��k
�Z+:��&��O<kc�T�'����<�J�j���g٬O`��l��k̼x2�J�#3g��y����D��#��3��!3��_#����p���+'������m����k5�sj5%g��36�Nֽ��Sxe����=��HČ� Ȇ����pd=9HFr�(�e��d���x�QW�6�0e�3v�&ϸ��Q��}�i�����qSI��'��e��������R��9��nfo���wI������6�9��|۵� rz��UJ>i$i;!!C�c`	F$�a� �Z��P)��Z��7�{�m��ރ}�T�覈ih�BF��r7����FF½C��]���j�(�|J��� Y�%Dk�)�u�Hp��.�b���T%5~���/�=cɗOT���).=�cJ*L;kZ]F1��O�b�aRkb���VS��8f�!��vM�{����C��jL��������ș�?��S%�0���/�ۺ�E��r�>�4����s9�R�E�|b^�|t���؅�O���r�h��mt7�N�I�])Y%��tM�t�h�����A�@Q޲�3عx$5I����㸬������5�7ym��{�w�B~n5��l�u�о�{i�=��^i^��%Do��S�<���(��#�#7]�"�O�������HB'=��#�b떱���}�����y�s~�0U�����X�S񦀚���`ЪGn�W��
HC����!{J�b!�a/ֱ�ۓҨ*��l�>ci��~�v��I�����G,�j|�t��%g�A��q�=<F^JR�	 ���f4:��SZ+vY��	?�����y��=�Pbx(E(�{{Gk\j�^J�-�^�q�j��؜k
ř�����������s��]V#:d.�|"�^jF�b	�[�CM�w���V�o�6�����~u��|%�P^� Y/���F��j�#��*@RK����-�	�9�cJR
s�e�����x�/�ևB�4�� ���:v>�B@���T
:=��|��v뉾p ŏ�M��L�$�c���|b�q�N��-�3L/���r����l��l��*���9�:���(��r��"��v�4�C�U
TTYah��*?J�Q���X݇��L�q��P��D��ϗ�&�C%)��q4{��� {����Q��{u����x��Y'������U��>2~�����I��>b�3�y��F�Ig<o�gѺ����I�$�ʥ'���6�+�o�2�M�;0x����js�ڼ���׫2P�zb�`wy��HޖՅN��4 yz=�R<��>:<��"�I�((�A�O�� �y%J��Ş��(���5����y�Qy��zP�r(q*� (�vQ��C��?S������׆4���u�=���|����7��0oJ�"�O�N���z`�V�"��~w��k����� ���ާ�[JB:E��K�;��AZ�\J��^B:W�ARR��᫟���g�;w��{�3w�L�~�G�6�d�0̽8�䄉ls/o�݌�щ���R.!J�������ߟ��|>Jg��I���>�1��;���S�A]s+I��Zj��w��EGJ����O��C��`w��Ż5Cx~��������Ѳ���!�>�ap�=�u@)yQ�H0��|� �'(��/���U\�]��l�R���$���u�gzd1����(UٜjGK;`E[����
��Sb̵n�x��C�:l���r�Ap0�����5!�.��wN��a>��w�F18���w��#�ﺑ������@YM��'/����[\thQ���_�C�̖�ЖZU<0+қ�-��K{�A�lѬu�p�5A��[қ7��2�n��犒g�~�� UW���I{+���@��C�-��&ذ�e�g��lXC�#�&Zһ���*�Q��,��.>聫:x�t��z\-��h~8d�v�X��?7�/�!~xJ�4���GB�a�6�6N-(^�xAٕ�w���+*m�OXk���=B���YO�;Q/z:���䪉+u�3�գ� ����Ib@�_�3��t2.�N/�4Et���"h�s��d�"F @p�����x]�L���{�P�`}$
6J�݊��,�՝��H����q�3�Ц������"fʦ� ��\#&(}v�7gMS��'v�Sy�1򫅬��׋E��S����=�m�hR�W���������`LlI��C�z�:�R�c.��ܾY«����4|�5���P#l�_��ϛ��
�ez��Ɲ�λ�C�*��tG��l�7:M-ED 0�m���V?�n������RԳ2Z��DM|�ڲ~p�w@󬂿5K_%��
�v��[���l	��륏&㗉ۤ�?�4?B��AA[��熑���ij=�\A'�,�@����г ^i��)���s��aĨ��.�j�^�p�u�mL�.�Xs�o(>����ꅺM��i�R�z\Q��|^���f�9�usj��\Mo���/:[Z���p��i���]��-�Shp�x3��'AX��~8�ٞ,١Fp]�L�����	�I���;'tY�~� ;T"�:��ᵷ!}`6�ou��j���$yo�e�wY�6R_Q.����?lm:���]��{5�t�A�Y[K�[���?m-��ӣ�-��ӏ�R[H�νg�^k%��-bF%����"AG��mfڊ���h��r��	3�+8u'f7�^�;�ß�1T�$��\@��jE����&�[��H�rI�mv�\Ǽ�̚(���z�t�̮L��=X����䀙,,��sk�Z��eX��Z�L 3ʖ	��{g�r;� U�J ����ٱ�,CL$ִ4��z���[E�D���{f�T,��%����\�+��J{�>+�����XA�QO�����~�)g��k�\�ԙ�%O��aoY��IvTAԕ��7y�.E��8�4��힪Źn~�w�p6�|�8%vk�6vG9E�#�}�}S�]�&U�3�u����&d{ӆ�m$�r�x��
��L�rj_eā��Y����M����D/�媃/4��$.����QU�Mp���:2O�q�E�np������"����Ill�=�@!����xrlXw�Oі�h��q�q@�������+�7�ao">Yp�-Mj~�I���I�u�e�%QFf�9VMQ��ޒw�Ô��=���|�M �@�R��Fo��:vN�7p�$�E�&���De9Lz�\�W�0��jS��R�r�+ûT��让��}~ؤ�� }� i��F�� �E��*D�*8�SY*u9&�y��g`�(���v�>sD�u��F���̖a\-��<+���0!֔&5N��J�.�OpV@� ��{ѝ�������(@�b�E1$�S�tvw��E���_~m���㇟?�}F�������{Zs��wK�Zd�����D��|x��[�B�Ҵl�D�Z\�>�E���
R��!�-��Y�K�v6�W����*��xR#��_��3}�.T�͏h�-1v�B�ٶH���O��|^gɺ/�r���ۡ�(������?�C]�䠆�N�
^R�uۤ��6�A�wn/�R�w�'�{#u��"�~"�s�f������FrD~��nϨ�V��W��g7�Ҧ�?�-#���UV�$��(j�eR�Q�ܻ���O*v��T��W%5���es7�&�.�0���Eu��n��6v��q/�Q���9뼛\��/�OO�F�^�t��A�=w�|�S���x,�n��K���~������3J����^��	�d���ۉ;���,�μ?���8)�#ϬV�:(dƃ9�'�dES�V���h��"Gܒ���S,�1��*[��]@ĵƎ��ך��  b=j�S����fe<1�N�S��i�����@���q3$���p���^ȖQ�1nMNL�`ηc��C_-�5@�S�ە�W�1�UL���~���*�������S&��;Eցl�5����W��U���Y$A6y$�R[c�Y�0Jqa��t�����,qɂ���}�ܸ��sV� �ɦ�6����;P����+�=[^i8�{d���v!��8�s�SAV�z��4��a��~$����-�7�����:��Ø�<o���6�����NH�}ElG�i�쎑(�#����-sr��`s��]e�֬���p��Œ�u��zAq~Q���9����b�ou�`_�s�=fd,cJ$
����!������R~��f�`�1���m�A�$9\�ޝGW���|3����2W� W_w=A`�{WzKQ;�B�B��~����7V�[)�l����j��~��#�Mir
�&�o�K�����~K���PG������5{�%	#Y�$�Ӄ��v��3~X�B� �w�(��wsTbO(�T)�|7���z��p�|9���4 и;������o�7V����V���e��"͑�x�K�u�ݔ��Y�_1Q��)�!}8��f"F��vl�HG)e���Z�[����(Ã���0�Y	���Ir������(o{�ˈ� ���X:��?��[|���7s��$���Q��n�Pd��I�]T���I�2��F�|	�M��,��@���:���������[q��x[�I	��i�/v����'<5݆�Z?i�m��Ct�.:�s�Gfa$��rtt���ywSD��H6)�Z���]N���D��������Q)�8�Ǯ�c�sb�q��d���;|ۇ�z�Km	.���D}�}�%�V��`��r8�f��$j����PO���h��q#��MK  �啁�l>�ӆ�C��|�XOU�us����w]�ma*}��2�ژ�E-�G���݅ٚ��Y�t�=��:���y��J�R)n��=vp���n��?>��|��1{d�����$~��q�3O���Kmd��uq�+|�&�4:������jiqk���uKH�yW��h%�0x�hYBq��N����f�n��>�9��_��,�,���?��o�P΂NMn1��9Ճ,�;}�\�"��@bp�����\ܗ�^���˶�8K5���|0��M֞��	�������pr(K和<BGh�q�(5Q�YCd~a�]�,�ŀ���}��g� � #O�C~�t��=!���/������<�=�E�: p��|���Q���6>\��78����lU����IJ�#����Y��"�-<T��f�L8d���L��ĉ�;��>0��e�啛��Iշ_ߕ�m����$�"�$��Y���ei���<ώg=Pl'A�g�Y.�U4m4���#$N�K��7W�W�e�x������چM��;c�HsgKb.�Y�6���.��f�� 1����OPr�]�0ֹXRm��IGmRŎǞ�5�D���1�-[;Ǧa���t�A�[�{�t�8�w��\�I����P��HM��d�o�Ţ+W��&Vm#�`WgK�JY��q�Þ����oT5���0�r(3y��Qlv�R��m�?8�߮�<�������5e�������M�+���U�6�D|���s�� [��t��˫���,n���V���Dx�73�W���Z��T�:�it��}O����3��ч�v~_]����wC$K�1��� �����V-RJ�zԋ���p���2��`�/V^��x��.�
{-�Z0�;L?�!0���ɼ5�ϪȈ�WVb��(���gu:En`�
�_>���A����pD�ArFy����<+_X0�h&ה��͇RT��/^Gm���{�]rr���*b����"M��wD�G��/U��6������6{�C% iMJ_���@�i����C��j���ݗ������ڦ�����ܻf��ψ%�0]W����5ިt��X�uK\��۶�����%�JYW�A�E��[N�W�� �pǦ�_k��o�۩�/��'=Ā1�Α>�t�?���F�0�{�x��9٥Ƈ���~7֊���`31����z}Y�R=�������9�ʴo9(9~x��Z�ꝲ�~W���9B(ӹx���Y�� �X�пYt�tAn!�m�����"µ�E�4m�0A��ō�f�^gY�/��za˒m���Z��a��{5�hdoEt�˖�W*��n:Y����8�]j��ݥ,�������c��0�*Bpӭ��?uY�m+ 'dϥ :s�q�f���(���!�qC��;�V��9����.(�)�[�E����..���>��;���~�|[�9b,qs��/�W6��n��u!\k������h�9���^'B�m����t��W�TN����c�>�cE��[��h/e}Y�ɋ5-Dƽ"�.�w�-r�~���ο�;��N�����uV�u�W.Ew�/��$��� s�TR���F7I���ħ�8*�*��>�fi�j�O/��bq����]�~o���n?��~ޑ��j��=�s�U����΄�>~����y�~�>a!Y٦DOǏ�ebP�VZlu)u�v�/'M���~h]�J �"y�(� d��u^b�*����%O�+�o"�)j����ƃ&�J��|e��j��zL����.H0�NVZ'V�,FV<�*-�}��%��¾XҔw�(��n�$+��,@�;�o Aʒ�0!�Y��e -;F�%�r�e�v��p �x�}�G��>�=�t�$�Bm�����Q��g88f1!wF���E��@cI�7��$L	�c�,G�(.2U��JK�}�&[�y뭊�bF�,�=����ieT���\�n��K�+�����=���1�;�w&A�K�ʢ�d�ϼ+�y˛�q�5�l�{{X|.���=���N�C���?������9�O�ؘ��F��P�,�1m�H���7|C��'���������� ���Rk ��*~-���r�.�	/������E�z������J��k��)Gf\p��m�s7�T��?l9U�v���Mj��iB[R�(�KX)~���J̒���7�g����/�i�۰i�	��&+�q۩�]nD��|a�<>�5�m�"��J�����)��#�Yvt}�a�,��1_����RN�$�Bc�JiRO�w��R�%�^)� �˥+§U��X�
�a���_����n�\~m�wkV��if$�h���G��J�w�y
����x�lY��ُ3�P4�4����p�}鶑���kv��B/�Z�rs�[�nM5���<-�Z�U$���Z
a��Qέ�DB=�&�ߒ��Z�7��P��d�9V��R�T�bM�T<�Z�%Z~���lt���BNZ�@o���A�.�n��	I�|l
��!�j���f��j�dz	�gzg�˟l3.�OT���@�?�gL��X�eL/'҅b�_m6�a���$Sg��U�l�铝�8�֠snΤ��a��\����UA�(�6��ɀ�]��/G��"��ޛc[4�z���w�)�@���&-N��g�n9�=;󠨲C�@e�b�R��:���d$����!��BD6z�ұ���{����U��n��ˮ�;.s��X�ZIϵ�<���3ܘ�П���d^��79gNC% c��j�QD���`,)�5S�-  ;�hˆna���n�?�x76��5�j�+��@���^���(�JO'nzD|h�Q��Ӈ���XE9����n�Bt̮/Ҩ����ο���+'�Q`@�Aސ�n��{����.j�x��F��
�77F����.>�+��KzC+�y�=렶�cf��Z ����0�����'��9!}u�SA�W�9QeT�QrJ��Tz�	^r�$�՝+.pt�5�����FP�f���Xb�Nm��4<���k]@t5s?ѴBxn�i�o�C�OoȾ���/ G��.��Im��/L����B��Ӝ���(ݛG�j�B���J	�qV�qq��ţC�cf"@"����?�����g=+��Z �f���ݱ;��|��fuU=�oٷkya��DWZgT��jFz��_�O0��R���:u�)�#Д_Q��2�ʛ��Ķ� BٕU�v�k��,Mɤ�+t���� �G'z������!��-GF�e�׊^��mf*��h�D�Q윂W�y�-�2��$u��z^�pf�R7գ�/N�I���-M����f�/�@�f�%���;��O�&��ZZ7}�/ݪ�y�;ͬ��=��1#���nt���􅢚�up'��/��+�e��:�v[l�L�<�н�;�}l�{�R�JTݚ7lWNnX�uv;�3��kV�kٽ���_ui vϖ?��M�A�QX0ʂ����	�F�@8|����A+���-tT��1^��
��+6:���_��]i���vj�3���}��W��@��D��2���k�Hb��+�w�O�EN���>��[u�+�T�B�
�k��,`0b?¾�Q��yQ�+ܭ���2�t�΂�x�Ғ�Fg�Y�h<Q� [�+��#���+d��\H/<il�_e�M��*zWe��%M��Y���Qc:�K�y�� �A�A�i-���=�ԋ���T�L�C�2u!hr`���{��Z}6@��*#n��;ԭ�&Z��=�t��l�4�+m�}�FD�R����<�X�Sv ��ݨ�:K��O��]�/�	���M�n��_�0��t��z{�����<td��<�}s�ПPP��u�\f#T��c�P�^��w!޺�_�y՜z�d��������>�c�L2{�V5��5�$(���gL/ �Q�)�𬧋w��1 T�5�r���-���]h�+�0@���Ш+d!]����=���*"��6]�~_�O��7�ܝ*����ZRZ�Q�W\�̞������J��7�����[8M�B��JE�A�G�C���F�é��Ǘjxtkw���_��f�ߕ{ƾ�_�U�w	s������.eu�����4�3�q�fO�����S@jI`�!{�^o���ݜ��vN���h���;��4�KCg�R���)�TT�o��(U"h� 
��Ӳ��|��s=��x*�i2�ֹͫ��4�]��뺯�W.B�H?���o4|��m��F��q-���Q`�������&� $E��'β�^7�֥d�:��G��ܹߢ�2Ćy�Tg9g��c����~r0;�}_#W��q�����ٱ�W}�x9E��3�d��l�^��j$-��� Ice(�;��}vi�=ª��4�:�(��"f���7]�eqW�B��Rth�a=U8A����4.�������ѻl�o�ed�|����m7�<����J&��)',����.��CM�uz��=�a�6�������	���L�/#;���rP|x˷�j�׻���O�O���v�hl��0���+fNbi�
�|ۆ�m�z���|�9��KXY��ʾT�2����g����?��/[��"�;j�-G�j �)I�� G��:�
�rMG���Q{�m���uko���$'���\ʷ��-/��~W*y���j�?ON#�m��J)���7�\��6�|)��[z��i> hoz����-��s<�)��M�Y7���׵�������,���~\�^�FG4���� b�yX#n�ͧ�~�(nja���}��y��b�3�ҹ7+���ڥ����"�a�w�#�xd�V�����̙�I����ù�<�-m����{#� ��~��	��\��@���"� �mi�:iS�F!���K���I-�o��4��L��x����$0+�s��70ɀ�;y�g���8�<��q�r�o�J?-��c`$?���00�~Qh8������w�w�1��Ol�� W�׳�t9�3z�7GB��]���L��=�b�=b^KU"	O��^�)��"c4�#n���f�4��a�%9���_���^���3˳��0��2]6��L:�݁���lt�tw��߇��;h�����x�/$VA�g�瑳�<Y95�g�/�+l~G�^�cz�H��������z|MxM _�K
C
�fUXF�j��jR�/��&�l�@��<*�#��>q�P��]��)�_B�#��B��|�~L���|xoa2�Y^���9�c�� �^ sd-�W
-�e)ܗe���΋�A�8M��9e�0� "
�����Q2Y�V�z �)<\
�U������@�x�����ͤ
l��s�D�7ν�x��
}�S�}x�T.#Y�@��n��0|���Ī������o�c�ૄ�w��i��D��
�@��X�5y�����r��q��W�J5`�(z�;i��]����Q,��0��Q����XLda���zk�{a����j���\mdl�=Q,�h�Tj`�d%p{i&t�)�+'7.��
�� K��=_ߵ�	3f�3��n+5�c���<��� �l�ܛ�>��7�:�l�œ>O����׼�`4M�>�N�X6�U�z��ź�a1���ibs@ڪ�}��}L�^�y��K$�N����ȯ��pd������b����s��R[*+x~7����r�iT�1
0[\���+�,�=�X)����f��Z�,l��0H����gx�ޝ����TO��+�B��?�z��a���o�1O"�lX$/&=˷T�K�B_�z2���D ���%�x;]����tc�]	��m�o�\R3�z�@�\�_��YfO��[P�@�������[��~y;�`8��z{�=/�0��̥ƘÜZ�6u�@P��|l��s����4_*.�hf ^��׻3a���e�s-H~�"�ԫ���ܨ��<������'�O6�M
���	��ZY��
��)��n�gg����VX<�x�xP� �Ue�O/���v�����H ;3�\���l2�мa�jv�Ώx�Z��m�� �����cI�q۹P�4�+��T�~4R�����>���Ď��c�K=��@��V|:L&v���{�_��/C�,ڕ�AV�(���V'�ºl�~%���5�d�#'����?�����}'Ymɘm����N2&��5���N�9��r�Z�K�Y���嘞\r����^���&�U�L*{�1�h0� �z�PX�w�f�PR�L��Ԥa�\����x��T�$�F���{��j����=a��� d#Z��ƨFI�B�y��u6��`�q��*ԞV��L㹔:�A{��A��B��($am������ο��m�`��+y��*W2S����gk�s ��Ԙǋ�$ӫ��5N%~����U��8͢�kI�kT!7�^!.�{^+���s� a���*G�e��Q�F'�Õr�ob���'I��o}�KF�r��<���|Zz-����	�$�+_B�n����W�qT'���LK6��k�T�-�K��g˛�N截0�j����rk�x��:N�]���h-�i�/f��{���߶��ּU�gO��ߣ[�� ��md��-�V��9�=��s��5��.�UU�� ��:���1��ߠ�
�E�.wn����(�Τ��/�>��Oe%�+��s"��N2�=cQ�{v�S�5�X��9�o>�<×��b��ͽ�h�b��ٻ�L�d�dک�ﵟ��eW|����pq-6�-���f[���z�`j���M���W�d"�9H��` �����8���@�����Df�X)���r6�.-oEf������������W�*�����W听�c��}�1z�o��"vv�8PB���/��E�7��M$��0a�����y�}�*��˭K����[Z �f�.wk���k>�^>�'��b��bF����a��o�ܰY���ڄ�7��3���O�G~zȍ�;���{ߍXf��w��d���&w��_E��y�#��.-�3�v1v���'��?��R��^������=W"�t�M���4���޳�\{��{I�ѱ���`�$BCpV��?���(nNԘf�ςph����[^ߔ�ڦ��Xj[c;{$ǹ���C���xs�Iz�K<����K� a���'�P������_�i��)��	Clz'fl��g?�XB��*�r���֮K$�?<`�g��� ��o�4k�@%%���E���?T7�g�q�i����0/@~�~dl}� TFY�@.� �|6���dD�T;"��نF(h�BV�E��}�����:1�_'ؿ�i��� ����3E`�'�����J�� �h�ʯ�!0�GG�g�b��+�x��_��Q�H�RJqɈcA_�C��<���U���!�eq���z��tr�h/���E�$>j�!���#�
�\A�ı�&�e;@��r�^���{��U��`s��@5�Ѵ��[�:�Q�� G~�l�)g�<��עE��q~o}s��������ży�eH)yE�7�z2�j}<�R	+���f�KJ�|���A{�����9<��~��Y6����w�9��#*�$|R�=�����,�䐴��To��Ċ�\�� !'� +!!O�n����rpg|���� ��3ns���h/yOA�9������o�{�"x?>\�|�zP�2�����C�֘�[�;�l6�P�=C���;�,>��}����@�Y���gEB��Т�(Ur2���A��f�	�.#	�8�^�����iE<d�|�?0�l)��Z>��f�$�!�K���أd�EV�;��E��Pr�<�!4�&k:�5f�BO�VP_��SDx=���d�^�\^c���A2��F��<&�L=|&�y�H���>iYӫ�T�d���zU�T�Ppܫ<a�:\N>/��Oi�=��Q�;�W`��[F��>��Z(X?'8�J��K�0�5�$�;���F2j,|$�B6����%��Eϡ.p�g�L{F|HH��"��g�Z��<N�>��CK�����9��+"�G4����5��T$����|?W��W=<�J�w��:0��x�P�he]�t��V�v����)m�?A8�h��{MX��k��p���mU����l���o�Z��ɗ9jy�a��w�5����r����y+�{M��J=�m�rɚϨ�6Df��g��o�
� P�^z�iBt'�e^Z+�F�c�.��NS+l�����I^	S#i�`Lhg�#�D})C��\m:X�I��p�WX�k;[+�R�N��,!.�M�����k���m���/��Fs��pE�}��U2��ρ���N,Q�DR�`Q?Ǡ&Ġ&G�BM�3����+M�#Ɨ,͐"��e�q�MlC��?Ϡ�j�0��m�`�WIc�5`�w�L<2S5���,ẉ��\D�%-��q��y�t�q���a`f�A���R�6��D�`m����+��̊ݱ�Ho�t�&)R/%K�eX�UvV�K4��R�$�:$u (7�ٶk�7�<<�TQ�C�E��r�CƲ�O�������/�܀{���Y��E�vYY�	�2�
�D)łT�<��ӛ�9>��#�Uӂ9H��<1��>dGr�DdBxo�Q#����]&��4�	DCK�#X�J�e��r���e:32�J�.f���]����
s~��:�Lш�j�t��p1;R)?�H�v��8xШ����B�r�@�|�-O� ���hy�o�ZU���Fkޑ�>���.�,a����@�52>r,��x�j�u����<^�e->�h�~d�5Z'ʈ��2{jD��K�0����3F�9Xpq��"m"K2n�f�E<�~�=v����8Z,O�@��3�#_F�Yy�Xs���[`�GE2��HI�����W�$���K4�Ħ%{�E��Ȟ���O�qr�uW��I�z6�M"�{������g�TTU<CE���Nŉ�!��,�X4(��w��H-���
�{�����ԕ��Q3�����܊i��+��;@�RR��}�ȮN��p�|o�J�3�.り�8���Ꞿ������w-���e��H�צ�cy
Zcy�yڥ����S
��K���M��dM�e�o��$l������Fb��Ipp�"Xa�?���FX����\�&�
p$����DGWYQ�eF2�r��as��%��x�vm��-s.�2����WɹP�P(����&�s-}l%�Qt8��3;?�w��ju�7���O�}���Y�d����B�ޱ��|J�)��գj"?�w��}ٔ�Y�*Sx�0-���4cЇ���$:0JJi��}���d_�L�7&U�*�zR[?��%Q�z���)IS�QF�rd��Q�3�.���b�;̇a�}f�H��}���2������&T-2}���M�	�O�x�ae�A�j|�ZϚDNe�ў�M��1���;�o���}���"=�o���T��Ik?S|_X��bj⯲`��1ޏ��Y��%��/QTS2,\%!E(r�����k]8z���?��b���A���@B1�,!=;z-������bP�k=���'z�)�XE)�GaI�����`wJ3���?IZ�|u2F��9l�m(�0�u§q���>�j�S��B�S��|}<�ۼ�J�>��HW	�~�=��M(R�����C�X܎��f�
>u�&�C$�i�6�����}�8��1�1�/�w�bʤ
�5�����X>T�p������_cfXE�#�nD��A�^v�k�n�;F//&����r���y�Y��g���>5`	n�}S2�ǵh�!Uևy(��!��s����*���޶~�'��Ȇc(5J������?72�P�-RkRrZ)**��GןJB��EG\����U���6S�-)����/�Z�1Xgy�o�"?�E���Ǚ�x64Y_�أk��xn��q[����|�m���������<�s-�U���.s8�B��tn��U�;���S%4�X|D�i�!��lZ�o͢R��e���Z�"n�P�MY?l&�gvy9�c9|zR�%OJ�K��Uj�����D/�g�F�� �ǟ��*Ԟw��.s��?�lVcK��za��J�,����a���zT%^�)@�\<�e_2��K��ss�|6*gB��
��r������eܡ؝#���x�ҙ@f�n�	�5ْ�ּQ��5�a��<v7�,I-0�� Lz���XM�}�%
\�jx�d�.&x2���xK~ǵ�t�q�S1���*ӧ�Zf�����b��%�Ů"��S�����	)Qotz	J~��O���_�
���:����T~�5�P>e� ���=U�&Fu| Ak��q����ڛ�e�');>�)��⅝�5��(c��G1죠&Ĩ���bU4[4e^m�+����t���O&&�x���S���^����wz�mñѻi計?|.�m�n~�_/��ę��ei�Yߢ�����9߾�����+X�u���WUb5)7��T/������ޏ�q��
RR��r���_��68Ț�X{niP�����������f�U��Kiz&�$���%9�C�@�ώ�f�b鷡a���M�෈��LH���]5��b�8�G<�}�{9���&a��>G$�/;�0	�U�#Gj��Yѐ����d��4������
��� N��q�f��m%?|T��{N��x��c�C/!|	�|[�Y }�F�X����r���he���!�b�nL��`B�����$2��oU��Pq��p�����,I$���9Mq��=�
ō�P�S���p�nދ�6D����x0�� �h#$�.��`.]|F�z���Y8�T����2X�A��m8Z&����%�?D�_lW�X��)�=�i�� |�(���LW�an1�v	�-�`����"6�OL�=0G�ȇX9c"a(�KY%*��G'V|����C�����{P诽��f�\A�A�*�؁���D�q�ye��B�֭��q���gqdx���(CC)�z9��P�t�@�e��"H��#e�o�	aȗ�xT�"V	�@��G�%ܞ5��x�c��>y��������0��X�%��tt/xY�*�eĀ�B/��Ø`�?�_�"*%bQi�v�u!-��nYjL��
&%��/CM[3p��C&�s�vǩ=׳ͷG������b޿7��|I���f�㟸�)�5V�b1�]S��ߤ|w 3��C{|~A��Sc��8*�t.2����wD��j���eV����S5��ݤx�7�b��t�i?�sg�v'	�I������J�"����눸�m�5�p�����i�[�W�坘h������ġ[@͈�wfB�(п�I{KO�޵R	P���~֊�9��>!윭3�£:F�&�5��1�5�>�YQkJ��6.m��<�}����bn�;ҧiM$	�Z�P�Z����{3�Ġ��@&���4�	��ݥ��IL��ߩk=˘��`�i�t�K��p�F���"Σ��I����}���qY�c��ix�� �52J哽�*9s�1��v����S9���������@D�GJ��i*G�Mt�2�@|�"�d~��P�q�̼�,�d� ��>ݩ�t�NJi�]�I�=�C�2�s"7����!����H��[�1��)��a`ڮ2�rݗP\i���z�5�x^�(��O��P+��[}H��PRuNWc 
T��t������GE%|��l�t�\�p;KY
����(�t\d��y&AD q�U����v�vo\̾I�^���HO�"�Q��Y�Պ����I����+���=��*��B�ؤs9M���a+E�j�7�f�����'��N�|L��]��Ör��yS�.��>�̼��p�Hf�>�͋����L!�Yhs�TC�-o��9|ע��
���#���"j�a`�W���l��AJ��40�ƫIM%���e��K��%�(,k·2-�� B�d50�u����g�i��|�C$*��S�߱��ˀ�ع�U������,�/���R��Ѷ 6F
A8�~��N�B�>�.��;&Բ�4*�\i�:"��Z��$�zz�(�/S����g������?j/����:�F�A.�xF��Ux?R�n�_0^�)���}?�_y�d��Z�t#��a�LF.��푀ԯ�Ƚ�f��	�UXZ��b�B2 bD?%X��{��KF.{��?�^֒�Hpi��2�°1h����B�Pu�?y�M�����$:�NAx�؄1w�v����Y�w2�O3�q�h� ��7�g=�#C4���¥�ΦX���!��?r�L������UQ2O��0�xeY�G�Ѥ��+�_BLu4K�Tn��)����ڳ+�q��������f+@��aD0��? �����C��,QT�&l�����M�IwbL�D���5j����m�� 5��.�1�4�w�z�����|�R�۰R葊v�%&e�ǥ�S���7j�4�SS,̀�ؘ!�0�ad��V,�$;A��$F.�	�N8��a�H){U�qf^&(���e+ҭ�� ���|�53N}�U����]�M�lO�V����0���򪄘��	�l�EdE?c KBt�a��Sq>eL������?���q�����N����3^D�gb0����^����ɋ|�%I��lm�9t�n�K���A����_|��h�1�(d�Ep�3ؔp�ɼ��[�
���E1�����fCMC�����~X����Mo	��Uϗ�Ӌ�n�_W}�%	�LBKA�~0ܼ{"�ԏ�B�]���j�@`D�n|y��l�j��q�?��}��M�
���+�8���䄰2��Nl�k~�)�H�ҵO��"\�Z�;�:ޜ�p��(���6d�;0��L<,�i��ⳙ!)�|�ԙƂhG3��"��;Ͳ��?���>�;��%����Չ�g31	)ɌW��Q��>vj �~e5�.�"�
��ú�n��#t���T�0娏���ú��S�K�C@����%�����&U��j)οi��|��Y��Afo-Wz<�s����h;;H�l'xͷE����U==�M�E��n����}_��~ �kTΰae%%	5�&����L�׾j�V�����CB-b�}0\���9��>ϋP���:P�T�%�*,!j��tR�2#�Z�,qx�� ��i�M]�.�T�D9}�;g�(�KM�sq����]�aju|��OB�"��Z,!�"��/��F�� �F1 �X�!��ڹ �2 �y+�P���|�~�)�D�:���к^,d���.��/
W��C'�[{.�ך�A�}*;���8�dH}6��޸�%����]���?SH��8ZqL�$��?iҵ�̼O��A�R�$p�!��3��<Ք{C�t���iGk�q>��/���`�l��G����.�v�t�bAL;,��M1�L/���u#.�|t�Ykd��� h]]���Z v�+^�iD��J�R�Pr���� w�Ո���=���Y�>�=�Q�uw�`�Y��a�k�Y��>��b�4�#�@��Š���s��k����6�Qpv,�הt��M��[۾[�.�Id%���⤙��+{�=�S_���MJw�4��4HI7H��(��]�"�2t�t!�twH��5��;���[/k�Z�1s�>{?;�{��Gp�9U\�XX���M�ĤT|"�-�&��P�!��B&Uϒ�t����9eV�����P]�YDp��3B_��_-��C�DG·��Ԙ'���Y��@�ظ�cߴq���vh��J�H��ϰ���*3��.�I� �2'���*��+�����u$�����|	�uFw����Z����Y����w��D��_�^�3�3<J�|��#�yODI����0�z��������
ǽ�1=��[Jx=�������Q�^�t�!��j�*V#Z���w�ߢ�����ݡ`�)�������5�J���Dh{�77VX�M�m��փ��V��~$P" O�"� M��o`"r�c�;{k3#j+����&@G�GO����h���l��=:`�o�s���<eH}���f/8��%��`kP��7�D���7����Y��w6rE~*0/�u,����rg{�:oH���y��;�X]�\?�<�&��]g����D^�r�ouw�r"m��B�q�ɀ��Z��Aq"�:�k����[�e�LtÝ���̻�)B5T����|AC+���YHq����:24�56V����@�x�,��j������I-�~~��^+���c�?D�h��kϪ�<�x���X�ҦO�LD�Ժ��e�B0c�CR��|���7L�_8Y�&K8%�Z��A��c㙜	�
�'�Ar-`�	����<;f~9rú������?���2�@����.C��]��7/3��K���YR>�1�6=��:�[��c6]`D2�����h()b7��4� '�T~����?Z@��P���Ip���޲��<^T|�'4�x���"z(�A}�	�}T�LӴv3w�����`���2�o%�Pzg������՚���!�2�?*�=\@����~�caڛ�Wx�]���$͠�ú�S�/�f����W�\v��D�}��ێ�V� ��__�?]k�誥�l>�j�Ȝ����/�M!'��r�Eb>��W�%ф������p�-cw���R2d�I����j��^�ky�d�)��^�p_+b���BE��?r���y��$�]��.W��
Y��'�/cmiq,�;�����}��C��q5����D��t%*Y�gm@�����~է��� /4�R4q���s��a�~7j:֗ef=������k��%i'�ᵭ��8̕HZ�Pu��Ǘ���;מ����2��(�<��:t�?ls�>:�G��������hH���T�=z]�K(8�D[�c�*�i���k��H�w��g���8�-D��ރ�5\j7$Xh��fY�D�Z�Ÿǎ��/Ţr��1���a��/�ݩ��G,�q�Br���F�v�q'7�
��J�9��j U(�kz������^M�ѓ�y,H&��ꀛ#�T���8�x��S�3l�]�4���5q��0��B=u8#F��ف�i�76�ĭ�щ�)�Z/j��Q����S�Wې��;0gw>�j���8�l)M%�1h;�Ĩ���ox��kc���O^�̾��~�g>?�g�Ba\,��2��C����nj���h��}����{C�^%��:�*m�d�JI�	��[B:ʏ,�4�F3R���"�@�Tr�4q�P��x0S�.�GU�h�}A�ኌ�Xkb���]��^���{�oG��p��%?��G�D'�A�j�ה�4QZq�!Z��..�~;7W"��9������"�^�.��t�9�]�/�Z��B<���53K�	�Qxxp���Z��	�ߗTi��2���g�us�6��Gaԉ��C/����h�	H��7�T�u���Oo�m�.����I�B|���L<��_���r6D�#	�sKF��_��.^<N�|�:�sƣI���F�M���𯆣C����Up��4S��f��ܠ�����������!�;�Vaj4�<ȫJV�/Ya�o7'���?��]"'������@���P$��F���.��s����DX��4��i[.�;�G�y�Jv��@��������� ,#��2���͝/�g;{�5M��D��*�L\T�ݽ�n}���g�+�׊���/��{��~�	G*���D�ib'��Yb���=[[�/G�U^�%��Q���@�{I��ؽ�����P~���:�\����+�%�������i��eu�~��5�
8Ħ������f^����s��SW�W��w��X�%Yq��>�7?:��8ܙm�.� xߥ4�]�|w3�����?	�Exh�K��Ћ  �����B]�^W���դ��w]*	-���4 �m�����{̀N,�{����G���@�N���m����}_X����*�jSN�1��,��}�������Q�m�H��$]V3�ճ�8��<^O����tܗ`�t=>�M}��U����L�e�A�i���3��D����jU��T^�B��й�F�CQ���=|�7��ʃ���K��랺����n��_Y�]�"{�8���l�	c�P�;.b_uu��1]��&�d)��{-� �D�\�u�;�^���b�1^N)R3F>���'BHv�(��Y��s�[:���}��Æ���/����Q��\�$�hC�bo�����q��CϵAD���q���^�$�p�D��*�DX��ECL�2\�Op@�f~$W���1��I�_U�NS�ES��lW>1�~��t]��9 �s���P�{ ��Y����T�!Än�� *=Mj��+��1`0a�+%,f��]#)u
��AGAr6!�̝�`��3g��Iwa!$)��k��x���~��u���x��˔��1��� 5�s�A�^]^�e��!����f����J�����"�uW,�h�Qd�W�	@�����ҿ�n�R��x+Y��f�	?GQքJѧM��}�t})v����,�R��2/&VԱ��0�ZZ�'����G�x^�9>��c��|��¼�qvN�C[�dM���Qu�H:F�]���;�i�o��=�<��/���Y,�`b��i&ё�/q�gC�6�D��=M4����T���dm��o�I����v�>;/���%WͬX3���M\��|Ed�nLQ�;4X�ĳGGR7Ͱ��@���=YYK�{�)� ��u�`ͦ $ �kC�N���B�Њ�8f�B|�����i=ޜ���]�}q����؛��K�y�g����ZL6{�Sx��G$�2����V�:��<7п�I�+��뱐u�{��g�,n�(+A�$�R���.��L!5�?¥��rjҧ�a!':T �0��$�ͥ&��^h��6�;v������^���-�
�7��Y<��E����f`�i�:���|�y=���E��r��)�~+��xp���>�{J��_�!r��d���[��0{���d�2,�,��W��u�'�
z�u�u{�g,�B]�q������7+��V���Η0�h$AF'�\$
O�!��np5�|�M��6O�`�;��9^<CK�4s|�W(ɿ���7�N"ڽ��!�xAV"��7_�RB
8E�ذ���<�SF�TV���fl���M,�9&�{h���ŚyO�B�C�o�J�ޠ��z��?}R���1ߦ�;�٫7֌�>r�cq��$H�}�[�2�Z��۲��'Z���*:��^)$eDYA��4ee���j�V���/��������4A\E�C�$�u=��}��r�~��U�)g��,_�ρX���p��=�jsFW1�!0���<�V��s�:�0�)z����
/��*��'n[2/��o�U���pX{��D?�M�������5��Pwn����0$ M�Iy뢏�dI�ώs�;����I���Vӧj���m$s�����R�u��/j~��="���^z�X����Xk2�+nG"�a+�U���{�G��oCuzd���}-�q�	����OO)3[�%&�̇8:G�&c��~��T����
�����>�ޗĞ��6�k8�eP�\_�]�^=Ѥ��iA�.pC���r��n7�8����z-�����Vh:I��E@ ��-�i1��m^�Ԣ|W�.�D�#=����v
%��޽KZL�."YG��r�K�=g����N}���Ђq��ֵ��7bpJ��Gy��y�<7[��d�髍��Oy�?������ّʹ7�=h<�����9�n��B6#9�+��y�;�f*'�?��-��g=�cG�EX�D?{,��-�4^��lS����V��{�z�Bʌ���#�RA���0��0�?�!��{����[*F�I�2<{��}�;K�Ȓ���m��j�.��XD�5��˒m�FO��������U�8�8�".z��Mީ�ϟ�Hث�7�+��a��pn^9����N���xx5'w���@e�JE��r#���:�Xoyg�H�bb�W@V�}�Bbd������κ��2��Gl�r�>��}ƽY
��qs7O�4�Ք��y'��{���"���?�ڜ�u�_�,��Wc����x{bg����AN����>���K�-G�cq�Im�91*k3�ρ�ث_ک�e'H�	+������p�n�^�gd�uÕ�!�L�/���![w(*���g�<�S:$�����T#~��׆"�tEq�\]6����Z�&&���������� �n�����[$^��I���zK���\�[��՘H�w��55�wTz��u�@������s��<�g&'����dr��ipY��I��	������П��j�0 ��5 ^W�Oݫ��l�V=`��:B������ƨ��8X��c�L��x�⿮�i�J�S�I��/��c�g=�|�([Wf #s�:Qzj����5ir=��FVF���>p+����&q��qmZ���4��]�L/hE���y�"�B���A蘁� �S�ˬ:/pӸ����/�
sT�E����y>����o���'��}Z��tǎUmM#H*���sQ����/62�uڤ�߁��Jǳ�*2��fg=���;^ɀ%�z�4k-H1�~�EZc�Qvҙ�� {���yvf ��K���v$�/����J�_�'�U;�[Z��8����Bd�rh^��fR/Q�C?�ɽn��&ӫDC�r��^��tNW1�0�Hd�cY]rS����,c��V�>�Cv��i����j�W\9�[>c"�zFR���2�bH��k�����ɹ��}/=�O��(�zۙ����{�?9?�%�ŢgiVO.�"�vh~�\��^�oV�BM�^�5Cg�~��p�b@��&s��x��e����/�a$U�֫�$J!��oq�b��
̞�X��L�����;s O�oQ�5�R�z5�lZ�M��1��S����&lYn[9���h�O����.&�b:�f�ǯ�Bl|�);�����;g4
g�V&�Ū�" ���٢������ %>ߞ������=�yS�[JFuϾ��͸���3kf�Z�g�+u�x �����ƮT�CO���Iv��F�"���"B@KWm�gM����Te)���Ԭ�7�>�W��70T\9�����7�L�9;�Η�b�g�Gc��9��I���xv��|'���R`0�0��32 �v}�d?6��lVݧE�4�&�^��"�ҵQ�IĦ�'P�nHܟ� ��$D�(�a6U�c�O~��Fsv�����g�~��U�7#���@�?^���<��n��zw��|5�7��{[�\M駖��}�B#GiF�r˕�I��S̙6��&�ޭ麋�kS�9�ۃ�pu���I=�GG7H�+��f�+��U�0)֧�$բ?��-2:R�f�kl���}�I'�������;������	Z��r���zgv�y��;뙓�;�u���E^�(2�?q�<�1k�Ďh��c�Ѧ�	���Z��R �����Y,M9m*��/b��#2o��H_,K4�-�(��<�O拓g�`�D��!Tm��s�m��Ϳ��F��Շ�u�HV��m@�G�y�"�)2/��>�������PAc";ڻW�_G��~)�����n?D���Z�D/��������&���5�&�n�	�i;Q�M���(5�Lz/��\�|�u��m�Hg:�F�n��%�U@����4�AFL��C��z���f�F�r�/D1'h�^�P�i�t�C /"���"eq��j?U˽Ʉ)3�d�����R%�b�Yع���1��;�:����N霝ؗ��Q�������:bx_�*ߗo8R�xr�<�����|/�[}}��Ef5H1:p���~q�<-/b�!@@�gd���Rد=�Z���%܂�����J����RG�:�|c��tP��P���KX'�߲PBN�����JkQ|1�Wn�e9]]a��z�,O��@��*r�8pՕ�/k:��@�����N��jT�(�r>1�6fSI-v�����k0Oۿ6���f|k�X�:�[��^4`9�ޟ�u< �I�e��9����Z�gVF;�3>��\l�I�Q�1~��d�"��6�g���9���F�U`��u��t"��y�`�������qs!����;>9,_�כ�3����31!G�w���5�J�6-t����$xr!���*���d��.��L�n�F�x5Ɍ��a��$���فg�ź;:��u��� �M�w�i)�Ot��k/�[�a),�X<�0)�jY��_��|�k�΂]T�g���� ���=��,�_��������$W4�  ���F@yg�/��=�J�#vKJW���S�YO�-Ę������OM���]�"S��p�_J�zP��V]VF82��z.P^Q���O{��!�!1_�C������N�g�>�����]ϙ\��||�<���ꅎ_O���N>9���Y+h�l}���9T��49�F�˾g��L�-5�����e҇p��іE�Ж>�y&�ط����G<V�}��!�{]�9}]6�Vr�D=#LM�b�>ݦ�[7޾��n���m�l�	�\b�����B@��1d7;hvul��E�xܮŹ[��at�����N�� 9⯵VX�h�����&,�6�y
�k���}8Y�`��9h�L=��!Oǰ��?�%�����g^T���v� �ă� �ѳU ��Ŋm��-�����3�Q�Ga��9�$-�e�_�=G�Y�=���˧ҍ��̞��))[h�k�f�6?��s\��Y^gU�sh��ȃ�`�o����3�K���ݓ�,��n�� ]5��u�wbxnM �X��=d�����jM�x����즬��*�}�mx���2����d:���KB���B��_H�P?�#p��Q߶?��J?� �#�����6@ܾ��]`�]�O���W�ݍmΏ�����޶Ծ�?��=)c��m�G:.'���s����g\P��Pa��VrӾ�X��kԞek7�h5Ѯ�dCMw퇷�12���p�Φ��_��p���W�]'4�Y�}o]�����H�SC?�нxm���;�/p8�9�J��~�����u�n�%Һ��'1��ܚʂ%������[�P�U-�/q¡���bSدRJ��c�V���ƪ/H�D�uVCw40]^�eտyy�,��(2�H����� *1�Q���v�D����|W&K=��rL^@�ft�S��jU�뙦e���������S�E�����_�^qt�Z��0�6�Ǽ�u"^ta�d���aZ��b�+��eV�I�	�����%���E��?��x�e&�k�.̛�����it�aQ0q�b߉i���4�bX��9E@2���Yo<^�3�?@��{l��,l��%�������gn�Ռ.�	�܏Ė�����~):�#�Й,6R��Y���D�v�g��я��L�F	�آ!-�&���g\\_
�K�~��%z�h���E�Õ�/��+�˝,�}+��<��B�-��]@!{\�PuR�L:μ�������Y�xThWgX3�U97P�3�kc����K��_��WE�=���݆<�oO}}���HƁ/�n�ް�|��ߞ��̣�N��oX��/92M���77�t�/�?�4�}#�-�K����xQkaT\m������۷���1���k���͎=���{��,`����\v�X��.s������T6����w�}B�H~�����[�\��=B�� ��-������|y�\k��	.�
���x�鰐�qeڳ?�nU�u����6�'GO~�6H�����'����M�Z�ۻ)�����nة�r�����֤��n�H�y1O��*��Nͱ�#���k��_�,J>�!f��j�wn}����oN@s��7.$+��������_��=���Q����o{8b7m��w�C�AxA�|���մ�#!��2����]0�)��*��w�U�N*1���4.��H�9�+��psj����t�P�	��K���Mr�Ϻ^Z[���<~�.�����?�>�{���uQ�Ǚa1�<���>\��<�	Idt_��ޫ=R47��~������|CYA�^6{S��-r����:���B����<"K2�F��{o ��ʑu2�� �=����?#}���:�i����Չ�˯�:18s�s������S�6�s�:W��4:	Z����^���o/�iI3�� ��a7^�y�]v���x�T�[\��2�>�M:/ˠ7O
�2�#e�J��R��im�<�2���%wHg������p�6�����㇜���A�+Y7�N��cjN���͊]�A�K�L"6�����"�<�)��	8j��r[p�����NW�d��y>R�%>�9����K܂J��4d���Y5U��p%�ϣ���I���Rݬ����R��u�>������W�x���km���.M���W��Lv�"����C�8��BWͩ{Or�!z2�F���sa;��z�f�[���� ��n=r�_��PV.t��1�(����0Y�G�j��؄6�Z�]2��K�E��@�ڞRz[SB��1,* f�Z�E�<�#��n�e��"�ti�����e���,�ֱ�<�5~uws�t/�i\���xk��*��E�\�h�+4��l8h���L��qM��,1b�������Ce�#��ӹ����_�D�|�><%T4u������e���qqt���]ښ�]���ਹ�=�+=�w�&�t�������|�rH��܎�v��1���s3��m�����0Ul�����5_����D�f��YZNA�YG"����g�����M��&d
=����3B ��B�V:A׆lR�&1W���P�k%-�ZF�����C���g�+��a{���:���4Ep����+I�d��q�i8�{�5�j�XN����C��$��ꂇu *�VG��V�Y���`�\&�_W�/=$��!+(���K�r���&�X�	�����c��R���~4c�������"Vc��c*鞥��
[�j"� -T���f*Jϣ~�B��g��j�-]��~Ñ��]�,l q��Qs�0���x��#��|�PqK�H12'`�N��_�s,k���9��w,��2q�H:�=�)���Z��7dX��g��RӸ~=��<�a
���^NE�:&�^���Q9=l���r7�L�qMƧ�N��4�/��_���~�1n�(*/\qx
�d'�:�c&♡�J�<��� �ؓs���L��6�]��!��#;7��5���^���D2�S`	�k����~�Ǡ@��qջ�Oy��Q�,9�
�k�q�uO=�FN�>���w\T����z��x�$�j���_��mB�|�䇸�#	��i�(����Gk���1��aHUu��|H6�Q�P��ܜ���@�v�����2&�QBс ��$�*�7w�N2�{�*w�e�A��1%S{kw%dV{l6���%���hIձ��؋�A��ς��}�Z����ڠ"3;i��
��K�t�7����䉣�z��i{VZ'ԡChjƝm�l��C9�������gl<�%e*����N��6�ȮA���Z��wP?���A��[��1��	�<�q���ḛ��Ԝ���4 /�[�-���q����E�Si]Mt���+�e�H�cd��x��o�__rvЁ�/�/�̢w�~F��뉎p99B��v��}���Hf��Iq�v�N~��XL�@ҸG,PA�x�$��2�5�@�B�1fLj���.K��i�@�@�����;ӣ�Q���1��#{Ut B�7����7{���s�����T<���.^2�o�N�{8P�K����9����>�w�1u��R�M��M�nI�[�N�ה��?a�d�}��r��:ڧ�b�E&���Y
ZA�Ӹ����w�����Uq�~}U
�;qC��iOZ ��fN棊 �ر�~�����C�F��*#/r��['&���x��ZW�8��,������ �ν�Տ�泞T�p���Z��l�\���$@�I�X.
�K�e-c�5F���hԛ
�� f�9 �^�W��ڞ	J�A�g��Q�-r�ga� ���k���u�qS�EVРk����T�\r�$����$�11�?��)����~�C�*(����c<����P�`��Tq��B��gr\Ou��O�|��E�Xs�8O�q�B�y��5	/4�I.� xV�x���o[�Y�c�7�i�%rm~0$�`j�[�'��Iq߹v����P�ܓ1�t��#�Wߕ9��:id3�(C\c�����Y����2E��p��9"����\՝���P�pBͯ~�I��0R����Mhl�N-����������f{�Tk�i�y1�+���^^����8����B��|���L���<�x<א�Rؽ�J���oj�n�%K<L��S#\m)�ϓsH�Q���`X�28�{HLm�o�v��aw�lk]2]\kMT]A���I^��W�|��n��	��������1��f�r*�&	������Z2�tD��Rb�IN5�������d����>}�gگ{%�=�[ ���_�Z��4�&:T�^}+(�?.�$@��������_�i��B=�c~������(=Eb��!�-�<���)��i��g�b`��u��{T�E��#����]�ۖ�o�A��qcu�3V���D4��L���yQ���������m֌ ���iYYJ�=�����XJH̸�{aS���O�,Ȧ��"�Ux�7�����ѹ�s�`�5^�h���0��>�2��:&�z�|O��QFyͱ�0��豤�Lo|��1�L��>�"�ʿD�T(�u`�01g��e��T�0q 	�_�eP�&P��։v谞���ӥ'\v�:+0����� ڲ�2�s�J�r^��{��u+������O�e\q;��Q�/�pb^2�pm��`�!��l�t��"! =u)hz &���e⍴D��ג!~�R�L!�׫ut�\�,m�^�-����~߃f�\׮}�O�5��'�T'�I��cD��	�|X��NA�۷�|<�d��¶L {�M�f�"ʳ
wf�t�'ܱ̊;"��K{B�R��J��*�|r�Ǡ��muR" &�X^���u7���UIN�{R�]����J��?�n��s��
�O�m�@����qԄ�ŐY�����E�^z�Ex!`���s̑�6�T�2�hv"Y2��QBN�C�}�6��"��܄|.�H�Ӓ�b������{ۄ���\�oo�����O�5)�:��8��E��$Y�1������>!KX���欱m�5�E�aj~��ϓ��g�ea3MT��0��Ԍ /7��+B��� N/�_RL-+��YGS>����},N���_If�%�?�\#VN4����*����[)){/d{���aa�5����j���"��ɓ,"�q���g��jx��f\oSJ����!n���2���z�l&���1$��˕����\�w�\��1���d'��֝�JoJ����n��,�6�de)�yO��|h'y�08��#���N��[A9X�(�9�2�[�  ����"&��2d�g���){AX�g�ϋ}�ӊ^��+�'��.���L?_~}>�u�´3��J�8�n���i����=N�P����S���r|���ӘR����b�Z�+n�W>��l����"$nÊbS]���<喎6���-q4�H�aW�m7ܐ�g�E��Gc�DD��0/��|i�GW�:�S__^�go\�7��H�w(���+N�� ���&�ٞ�!I&Q�7�"?o"E�.E)�(��*Ðd����b d��$�	IQlQz�G=�<.OTD�2�B��t�k������X�Ġ�7U�7lj��~g��z�eځ⢩@��f���F_��}�E&�	#9���skN�Is�&t��)���M��bI�or5D�uJdcɔ��������vf�c蛼����J�?q�Tr���;D�q�"0�M# M�
ctLX�{�7r��PP���.�s7u"���h/ַ���"���ζ��|���������#��\�q��]N����#���`�h��$\~��wy���h�,z��K��+�����������R]������i��[*��e�����m����t5:&�pºl�	S�wߺ�a�U'�u��;���tb��w"��o�0�e�8�F4S�UdQܧ�y.�j�5�v�m���"[��.{@`ЌYg"�r㵡��z,*�l)��(]ٴ[Z�c{|k(WC�."Ӥ�x�N�Pܔ��`d21�u�_|eśG�K	����O+�#����\�eR$@�Gz>�k`hEI�e�S�D �Ҟ��4ʏ��A�ֽz�j�I?��id4.1c�ϩ�!��`'�ۈ;&��٪^������b����9�F�7����?oUL8ӿ��:����'��ʐ���{����B�%gS�t�-X~] ;֓(;����m�b��V����?>L��F�h�bN�ޟ"�;�D���!(��GLB���wh����6��S�6��=��'a<��;�J�n�qn���l���oٽ�gYrڬ����+s�7Η0p]X�^DK�b�OYB��L��hbyVxw��jU�W m���B�r��N�������.�5�*h7���p�Ԍ��̦��_��!�W7���D�%F���<��8H�Ř^��wd����$�F���gP�wC@_��>���>���+���g�z�a,?8�fn�C4���T��ɌQ�&��`�_k�N�caFZc���`��5H��d�C�dP7�t0��l��zRR�(IMȠ���bԒe<�}��e�x����y�)��k@�Cc� ebT�[(�-���Q����1�߸�s�_f��F�lmkL+$��
!I�U$�%?���9n��E�\~E���������u�{�
I
��}I��A#����@i���8.83��\%VP�;��(�[�=-��}ǥ������g%�C~�CP �ə��W_ߘ:���1�M;B�"��浲�������З���K);Ȝ �I�c�UR|1b������y)-�|6�#ʠ�����+Ln��u��z�M�<]78�"� c�;n����<{�fU�����iC�l�O�+9��A�2J����[���U澂2YD��٫��!��΂��({�8�Wf�
��In��L.wk������Qz�l�\�%���1���p�����{V��q�����0�AS�J����:=-��vo^�掐���J/�9
zƭ�5 Q��1��!"S���$��X���-����@z���ixu��y@�xF��HQ��f�9���i�����u��1��`J��ᩇr�O/�Kf�n��Hi{n�C�VQoA���{4���&{;�I��F�g�Q�- ��r=y�g��Ss�Xw�$z ���3���U���e9]bQP�i.�F"��X_���
F�\.@!t!#1��
�Hn=��T�&����z'v��u�����l?1u`�ġ'B��r���?��r7N�ag�DYy
!�XQP�� S�=��m�x������M�=;ǯ*n�A�O_�_?I�!9�T@I0��p�o+�(��VFp�KV|����f}p;�V)���U��饧�N��ۣ�Җ}�[�@��[~�K
mB��Dom��1�����pX��8�����ܩ]wgu�g0��y�1���¿r�=,욓7I�=��MҾ�@��E��Qb1p�߹yx�W?��d��&�7��m	�L6���|C���a���g9�������yJV[���$@u���M����
�M���@]R��q��rkg/�.�dKD�f�"�9{#蜢4Yad���x������V����M�L�X�i�����j�	O��f���4�����bq&��D>��0o,��;�O�� �j�ܘY�\�a�'��A�t��Z���3�}�wP��Rq^�i{P�P,��p0���F�}���vX�X��(����RS��չ��S�(,�9�������� g[�e��V������@S�h���ow��G�>���2f7_��>�X�;�$��t6�П-���=8��X�G/qf>��4L�l�|wB��#��ړƹ��e~�L�eC'�w�-,�M�?L�}�h׾;f��0���F�)�f��$�k�p�F���(���\����?�{q5j��k��턲T��$f`�P#���y�j���|��#� �*��4�������{���{��ʿ�'���U_񽏘ߤ?As;cۂ܍�=�"��|
j���|''�шZ�`�?��]m�m��Ȁl��vc�$l��8}�K���ٳW�/�<.�;�ڳ���W����U`� ;�����P�ُt��?�E�UJ��xY�V��	�{`Tb)��}*x�x��~:u���;GĨu���y�������U�O��Щ�P��.+Sjl���75 3z�D)]�ҀN߶�+O���2�T��b/s29V�W�T�9	�,�����4T������kF^\_��X�4���--=�S�b�����'6%>1�ք��|7�d&�L�$g��U2[�j ��P�����,��/SZ��"T������h�o�����YE��H��OJ�'y��'����}�=՛I>�z쩔щ�L
�Z��-�ў���`=|T�����vi�s7�*ݧ6,XCn�L�t��>��MO"������M�@�^�N���W�������@��3�>sђ�l�a]��:o"�>~����;���$�v�6	3����>؊�&g��=[�� �B@��Z�����3���}�,L���ѴM��D�K7��N�$Ҫ�����^3���g��t�a���-jӐU:SA�T�V9�p���
-|�,d���"#���jA
<���\��aGc��r�vW����2#�԰m�4v���{�o�9�3�L�􉐆���h'+XM��3F�'�|M9JQ
�6�07�������uyjƦ�7qO��;���6�,x�w���h7�S������}�>5��7�*[/�i[ �c��buq���38�[v	e��V�B�J��z���-��[Nh��2�]s}����6����CV�[����HA�t������ڕ�t*��ܽ��3rp��Vh5pX�Uޣ]
�"����q�a���'/����Dj`,җ6�>B��+�^p�ZCX��:�/Hi+,{�� G����n^_�]gbr�!���k{KPv�I� J��r��b�\�v(�N����_�~��=��:�� n��~�2>cם�����2.��=�9�%Tt��g��IH*�]��w��� \7Zwfޔ!���ܠ`��,�W�f��;�%���ƿ+��@�����S�b����]R�T&j������~5���?�l׎����Q'5qՐ(+ث��.���� ��.SR�h�=�v�J�ր��q$���Pa�z�=S�Q�>�O����]_���%D��3���p�6�w˄�y�O�v_ӮvQt��&���x%�qڧ��;��D��B����1^<���g��]WQ�o"�n�s'4�,��f�gʢ����C��g���׊i�)r���G"z�h҂�a�����9��l7��"�a�B�·����D<l>-�ZO�x�Ot��V��&},�(�s�̦�{�l���1�����)�HE5dp�^��y�N/���k�g�wyA�7N*OOe�<����Y��r��r}��_sQ��
��C
�C�.��ӋD:C�r�������|Tk����(	�:��r��UP�V����pY8:���3�����8g�ٽNH��5�ۼ�|��L#�dQa��&���{(��<^�f��]'�a%!]y���ϰ���	������-�S�w�����a9\���6��>x�	�����0~��E�{��*��0z�=Ì������̓�i��b��D.'/\آՖ�+���S��Ŏ�b�E�J[�~�O����&�wT�>���cR��,�8U��F'��3��op|X�����ZjP�u�>lVK�W��ꚹ,�&��Q��ͧ�NHv�[z,;m�Id�eao������&�a�p�Ĝ�LXn~^oKѫ,)W���!�_B�>x��Pݓ~^ +/̩�2�!~'�xu�|8�6f��ʎ�"/��	�Y����6��QU�S�WVF4�82?���԰�\ۀ�KM[ぶ7��>��t��g߁o9Y6�h˦rpj�B�8�iWE��� ��Rҥ��)!����݈4���Hw�!�A:!� �xo��{��χ�f��{�u��5�d��)�`<��������m�ý��q�3���J�Uk3͠��9�z��{joJ�C����ҵ��˜�y�=i9��,}���5�'��nWm1��\Ȓ F��tq�!)m�ǣ�(>�}���d�^~���_�1��4�����侸UfYb��s�t��ࡐl� ���iڕƏ[���qI�/f���U����^�����9����^%��j~�5�z���-��ⅆ�&�
Շ�˶8J��4�b2��ə�'3�6b�'�hB�H�*�ܳ
^Ֆ�6���ri�o_�'���V/|^���:-Ȍͩ�� ��XC&��қi�sd�V~�e!���tse! s�FI�}E_�K/`��x���{.��>����@�a?�{�a�wmo)3�p��U� ��Xk�����q�Q��O���e�	)7w������s�A�@*�}*T^�gn�X�R�V�zx����X>nJ���hb����iÌ9>��R�3pa!6$�/Kl���������v�]�!ۏk��x�fb�t��o5	�}n�e��%�{u<�DI�E.���Z?x��~�u\���v�Y��H��w:�����%���$w8@1�\7��xO�#�l������g��*���sx�SV|���O�����)G�z~�v%��=����w�M�+4��Ѹ�y�󸪖LN[)���_A/���IKO��rs���[���&�p64z�m�\5��A��M�� ��[���}k��CEw⭷�ɉ �/w�w�z-SdvBض��8Ɯy�����$ǯ��m�d	�80##�P�5�;�![��ȍ�I�����{�C�5�V|N�z��qZ���v�=�Z]6=8�3�DN(*��P�m��YP��ТI�$`<P����E+ɕɶxDs���/D+Z�s�E�i�DAE�R!E4,�u��x#��q�F�P�/�"m��# ���♫��^_K��6��u�޳��]��4����t��\J�f�@���Jy�=��!�0NRw����ֵ$Y��_�SLb�X�4}�U�F�5�C��4� ��H�h�S�K����2"�����̻!��bJMA�W�DR�X].ɥ��}~��G����udF�tJ�3�����o��ʂ�[g�M�l�r(jH��u�{���R��[�A�q����tK���Zq���L��"���^r|HNeR`n)i9���^[�rF8~�W3F���O@3��ϣz>�&���h�J�k�����{ڷ�7nc�^��S/�?� �1M�p/�+W:Vet�r�)�\�_����@]� �.HW��f
� Ɲ�4�h"&�JFP���X'�n�N.P��h��g�Q�)�0!��nX|��$� ����Y�yc��/ЙַK�I���u���7���d�����nQ@�]d��~A1,'�̓�[�6�*�)7�r84�<J'O��i�zw[|�-�T���'��։Z7����0}��3j��lzhY�:��d1ׁ�����H�)�~��YPJч����5��;E�?ۃ��g�CG��d+W�#�Z�j�ܭ�Xl�_�Y�(h����`lC$:=���lG���o�}r���O�`�%Sk�Sw���~�Iq����G}R���5U������7kR�i4�q>�g����2�Kk�I ɴ�-ݸ���,	3n ��t�+�1 )HU`��]�EV�#C���>�<�w����hl�.O\��h��̭���5��낦K?��n�Cz��v�F+�c�|�%l3�j!M��`m}�����rh{�	q������9��_��m�t�o��IB�{�h.Sgu���"c�����:9(y��C����ADco����Fd�?��EU�j��e�TS?���\�3��⊐>j���[�ނk%��J<Թ�]�6<���<��^���#�� ��Ô��~ߓʠ�*��j�$U�w�Iʥ����ir�CJ���g�h�+��b�ݣ������$�N�rV�c"jm1����8~�Q���I.|k\v��^8�����[+z����f�+x���!;2�PX#��~B�1V��P;"]~�ዦ��>;8G���L�wAq�*�)�
WU$3��ϐ�Mn_���Ck\�X�-���}'ᑆf�{������X~��E
�Oƥb)�K��(~d��P�����S�Ū�.56�\��/<�T��8�]��>����T�a\�5>�2����x*Χ#����91�97_���	ڒZ�����)0��M�+[�+eY��Lб9��d�����s?:���km�w�IY*�,����۞:�o����kk�+s(�8|��,m���]M`�ԉ����<0g�)o&�sm1�7�J�"K�S���!�6����E)���� �I�Ak`�1n�࠯�؈�_��	�3?�7)<џg2g�Q�]�����SHe֟��)U�>�f�(R�2��1ܷ
maLvűkdr��sy7k|�����ʇ�%��XN�R��!H��*��5�,��x_L<y�?÷h��-��4���D'#7$/��U '�_h��~�7�R��݁/�	������`���H[�j��b�	XZ4��<��%Ng����rA�=`�WEqt�֩H�)§�������d�uث�_�9h��!y����zq�zICC*[� �jgU�պ�n��&R�^ ��6S�o��e�є�;bg�S��x�L�?S��{G*��M�����D1��ڇ2���m��熪�ǩ�4B`�T��=/���K7�'���	�,���4b�kB�D-8��&>Ӯ��	z,r̄C�M�F��-eg�Ζ�ҧH"匦T>$&��ԅ�wSb:��Yh�)A����/�DU�,�u��SL����J�΋�=LYT��߂ZN�Zf���R$�&;��@3���*�Vt�Ow�cSV�=���*��ݳ�����붠J���	z���L�0�IF�\DR6�P��N&@,ж����p��|镥Q��c|�71��|�Z�'1�X�]v��HZ�>Py\܀��_/��a�a}lK)�v����G��h�:��ƄQ�4��ԧ������a�:wMJ�O�
���\����f�0�����\[��������v�A⩔}��|@�O>5��n�w9
��_{5����?F���k^���3���V,��sX-�h4#��d]O>�ի�m�~�Un�w�>����tTK���l;���D����'?6Dѯ
�h��@j�F4��x �*b�c���:�
E������P��	L!.��[K��`��%�a>>���>��aSX��t~�PB1��z��ka]A��Ok��A���\��6��N|ѵ�{�����8��$Q������Y �ΰ�39E����o��/W�#��
a�cE��x�b�s��X�ν�S��*mWoa��jg^rC�ئ#1qL%D�V?����U��n�^�W�S{A��C���;�-���|#+W�b����^�=�U��Xs��ۚ��4��J�`棧�N$���Q�fh��^oxBZ���l�ȼ�V�ү�*�����MN�#�a��ǀH~��>�y֮�'D����`����$5��q���h���X��+�_#H�?�z��M���a���sO�(m�$�&�sD���FtMr;��Z���N |�n'�&���yk��fCFA�E�篝�%��|E}�׿����e?���1P�3�<�K�f��k9h�!�kZ*�5G��t5Js&���z��_L�YY��4��ǐ�kME��kɗ��=,w�F7 ��͜]�b>z�����CNN�Dr��UP�9�X՝SD9	��wz���Z����Vw��,GAs����,F�SHNB�C4QGz&m�Te#�r��虥�jb�\�*m;֨M ����[�2�f�D�{�/�� :ֿN�wS����չt��O\]|��:��M��.�A6ҩ/,�p '�8�0H��g�ab7
�<�J"9�R�^��iF(�d��}�~$˔"p�	9=���,�r%��]��cc�?�<󜽄�ۄh������#C9�#�Vx��ި����[|{#��&/P�e���eΧS��^DK%xфP\�=��脰y�Chrۓֺ�����S��}HX]6��g��﵇f�C>F��#Oݱ�>�oH�6!H����v~wON![yQ-�%ͭ�"��G��|M�uBqyvp�up�p�up��q�Iqy�p��qxH���eE>�B�2Uԟl$n�a��Į� � //�+_�>Gn᠁�K	���}�2u2�Jz��X�2_��o����}�È�n�v�$�gz���S����+����t�#��,,�{���t���D�	�������ʷ����wH4�N3��5�2��{��c��U�����l�o�7498B�#���7T��D����ߤ'�8���?�(�[���D��nHD|_��S�~}*�c���#��d�LqYY��f�D���Qqq���OA�,�Y�X�XG�L���IUg9�6\\\,��I84<��}h����'bbF��y���!}���v ��G8^���׍GS;956��&&�Se%�����U+�Q�Ɔ	�,��S��� !
,	9u���i�͡��u�����ke)b1a���uD>������d��4S����/*JJPs�H��tӸ=�ub���,�À0_�qN4{�ѡ8���L��0""���i�0�!!!������F3�(Z+������do�B(2[e��;�(H�go����j4�"T�����F> �1��Jyx� �QWW��A# "�L��.������G߻�ߦӳ���V�a��^�03`�x�u�c�<�jf	��M[wmYsLJOGNFlZ�)�j;�g��g��n���K�NOO���C��R����_JF�?�2qr�)(�Ƽ{w.����MV돥��j�S[6����M����� ����א+���6r0�̾y>��ݹ�˦/y��=/�������lD�lD�+{�L=�\��L���WWWKK� ������
̊��hق�[�?o@B����1C���{�����H���S���	�~�ͭ�d����D���?����@���>:�����l���Jjk���݋L��fd� ̎p{��(|n ]��Va<:>>=��(r�Nkggw.���a��h@�f�{(�%���
�tD���F-aC)9�TOSP���������P��@u@@��o�ί_�p+}}r_?���瀃��ϥުz����i<�?N���!@ )���:y$�:Y��{����N�Xԍ%�g	ǩ��2
8f���y'q'	ӻ���x��?~��$H�W7�
{
AZ��pʖP��ǟn�~�������}C-�(Q���gسN���`�?������͵����!&ޟ�P��,\�x��7ر���h������*�������?[�R���:	B0���@�Bֲ`�
�V�����|ɘȦ�'��v_4�PQ�sKw��O��	�oC�*y�����R%���W��V�dÅQ�����OQ������/������1�cQ�o�\��c�����ƋKK�O��������7k����������	���Dм�ڳ�����L.�yް����@� �n���Ω��da��nx�+�����mGqv'4�0�ya3r,lH(}ښ�։/uőI�����D�c3���ve����O����=����YY�jb��o�S�������#�jo+���b�LSUؖ5�k�Ix�"���EK�V�v�E���|Bq���1*ro�k5C7]�=���{*m�x��@�oOw{Pك��8��U����;ǅ��ʃ�|zv�Bl�s�	B�^�@Z����ߌ�\��������z~2��� �}�
�.��m�}t�AȷVM5)����JN�ͣT����A��88W	\eD�l׭��QNZ;�3/o;Q9����ĮT����hVd�Ƚ�&�([)����O�.4MŚ*��v�Յ����5?ݎf3
?���v4�������}I��H5�3�������L1��_���a��Z"�� ��AQ��W.zy�Eʕ+@��8*�a�:��}�S���'+:Qk��8�B��2�d'�v���\7����4������[-z�%��Q��x9��z S-��U��J�jҠ%q6����j#7�����w��B��NO��4����wI\پOٶ��n�k2]ukV���ϭ��8`J[�p�y|%ߓ��a[�����6��g�b��UkF;���-z�+�W%�G��u����'19;�2��r/���@)�~Fp����_��C? Q�ld�
����)�BB	������X�˒J�1�5�h��r��3��K�`h�X��ٓ��뱕[�l.���0J�5ۏ
�|�M���b��WpŊH�g�>����z�Wl��W�c����\�H�UQ��Ǆ��﫣AWH$���/e|���O�2�N�����y^�=�k�s:��-���-\�W�.�R��sO��	���C�oa��m��Y�yģ�I����ȃL�O�d�*���Lr�C��w{�X�G���e�e_�f��^?�oU�S��8uf��_��A�*�g�$�G�=�Y�WW�(�b��_Q���b������]K�������5�����b"x�.��]��ֹ�L�'i�����%Hh�}���{?A�� �<�U�U� ��C�����m��$Yb�bq��.UQ�-���oj��\��m�;S��ۋ;c
1��Ggc�����ݢ�@�YX�O�;k�0�8o�{��j�%��b�;�	&?�������hێׯfr���ؖd�V��7C��AJ���ˣV*2��n��OJ̾�O����t�\�Ο��FJf���-&������s��Ժ�/#(�E8�;��N)#]vA��V��7j��bb���9[���̄o�	�/D)�nQ����/GF���&�b�+�p|_ufB!�����/��{jP����F�N��M�=��@
�JԵbi�<Tx8z��Ik$�LٌQތ-�W���I�O�.h�S:#s�VBt�*�Ga/و�)+so��G9������K�K�N�j�{�ߎ!1�6�$)o��B��&n�	�8��S2�ˬs,�;��,X�ɨ�9�{��.-�:݉�:KJ���|SO�y�oR#����w��k����x�i6�C�'̂��w�^�a�!�"v��G�L�ρAa��J�r�u�B!����m~۞�c��Qp�_,�E���Ͻ�T�ׇ��~��C�%��!�*�0/l	m=`o�L1���O����9���>U!���{�83r*�F��a��ª�1H�6�(���a��
��o�-����HT;�o1�v�]UJ5����~� L��?b ho]|{�D������ǭ�1k��"��>)5=�GR&/l�A���`m��P($��>���V�&CO�,1X����QJ
��ŴCd��k�\� ��I�EϹ|/v�r]�du5���uv����&䱒���pŒEArW�w��7�]uH��lël,�p��ת?�����иO��*�s4�a�S�	b-�߽Vlקd[�/+���듧�MND�rS��U���q�}~+����i6��Y��I���5邥�IX�4S�QAe�=Ŷ���U��@V���FDe�az��4��M��^�����/ì4#ף��IxY�7:Fi�.�1�є����
�7͚�$z���\�~�~��i�"|��j#��^!J��{V�<�>�z[dB­���l��m���i�0�,%F������f1d\4�"L���*ɳ�o�>�)�?h�ɉ�}=J�7��?��n����f���FC�f<϶��R��QNi�ӿ�P��Mv�9�:��f��;O��b���u�s���������������<O�T6��}�����+r��yn��oIDmi�bX����U@%��BڜB���Io3~b��TⱈM�UB�㶠�� ���zrq�5�̋�AJ.+��i�F�m���hx�)���ZXH�x��F��qAdȪ��Aӗ{�1��8{KǷ��*{��ᡢ�:0n���>�~�g75]�
R�"�H�����V��ʐԙԘQ��}�Dn���cE�E(;�Xo�&utO8�cC����g�pfW?�g��kT}ڋ���e�������vzT�~� "NF�-�;��:[���s8�}i7�2p��6�r�0�&r��Jo���9Y�ժ䜃6�V;���e��ɺ �?���ɰ���d�f{_t�\��v֏���]��B�o��	�aD��7�<64�^5/U���/AT����Q>��4�n�Q����so���{�۽�Y��yM�A�G�|

ٍQZ�9�p����+�������r�0�kĴ���k�����UZ2S��c�i�z�wuՖ��;Ǘ� �K�5DsgmZ������V��Z�1�Lg��q�§�Y=�ݵ���7�b�,�V�˶�6���
�5h2
��HȜ��`���m&�����¯:MWR��X���z[#��/u��>�F7�*b��L%*�Y��ȗ��K�Q;�3̹����c�]ow�mX��3=*�q���4��8�Z��Br��_������2B���	K*y��W���tH�vn�p�����lm�=-�t$�A�B��gF$��G-��)�˔M`�%�J�K��`�a���}Q�O_�;���`�/f�������X}9�&4��EP-�C^�T���d�]#�k�I9�y"�ft�k�ר	v�27�v�V�Vj��^��gaۖV��
���;��fM��k�Y�,ms-��;�GIԇҩ���_o��b��r"L�}UjX��?B�/MueԫMF%ۯ��V�sn!�w1���l���ĻC�X
���A�Zz?��r��J0ju.���}[$A�[��חV~t+��:��c�?��,aI~���N4Ϡ�� ���mB�v����	�&�)n�P:`zo� W�.��f�ȟ����C��=O�#%��sD������>.+h��R��(-5=�vろF���~��Z�N�����V�zx�K�]͛C�;
�M,��sn�U�}(e�i��]�;�}|���Qn�������{,���� Ij�!O~��3��v%ho���P�N(�1��lh��'wI�O(�?>TTE�m\�u�����n��⭫=ap�Hox�8��y�����oT�g�ˠ;b�w<n�q�=F�q��P�����&�:�;q��sU�;b��Z6c�ύ�OL�SG�}1�n�>M��=ȗTՈ�'�-y2#�w����ę�# Z��m0@�ӓ�6B-Æ]�D��gk���s =`&���x�u��K�����s�5��Q%�P�\�w1g�v�}�5H}���f��~� I����XU�|���l���wa�,�ka3������ۃ�	�J��C��ʮ,/���b���$'��ؕ�Ƴ���Q>��*�?��B-DL�����b�jͦ�H�)A��W=�/!�����|���H�=����F�ط<Uܳ$A�:8f��xWd<~�R;|�Y�6e5vy#�&c�� 2>"P�T9<�dus��~�s,,�HS���	���6��]$H��~��%j#�\{*]��2�}�������`�3�]���v5�f]̚�x��ڵ��\��跒���"OG�L�on�=t��Ơ�_ZJ�r1��XM�s�'4�N!�)��k��"T�MOt�ٕ7���
E��D�g��ť�O��ku��~�����0IqYu\6�\C�W`�69���6�k`����(���6�x�>�gћg���ލ�_�GFd���I�꩛���v.Ծ��xK�vUs�Z_�쩋�'^OL������'G2u Z"}^K����d�񽤛B��DTan{�C[����sɡ0U��wX˘H�w��Q��\	���#EV�2�j��d�}��7��;�_jti}���@Ŋ���l�>�z3�#@�#s\�5�4��@�?V��Q~Mh�/��`'��ۻo�!c�UQ_��K�x��dV��
u4Hs�|����S >$_ ����aYi�i1�+��P�{�Щϼ�E_۰N��T���l�]W��K�����|����h��������/j�v� U/ ^��嗀_���}(�v�|��;`
����t����(�v�<�r(f(�;�3&�,k��X�{J/v�����~|�!��G�9�-@���|1=6%�F�z=f0%�?(C�!u[3�+����+�Y��rH�>v�HB* b�����Z��`��w�]`�M�6^fKи����x�e��d\�?j;����
�F�����|���w�41^u�
��!4bi���q�n�e3	/`���.p����(�ȅ���)��5���Cwr��JS�y͓�� ��R�M[�쮠W�9�g��]��Vވ[?�_����&��-$u�g[��&Y+�����d���pm���"U-v��;�s�W�G��u�p����y�3%F��5Ty���o�Wh�WH�mcߦ�D�(_�4`P�¦u{��	�B��	t�I�8�LN����PQ��oJ*�zG�EX�yP~d�Xz�E��6 7�|}K_<i��Ms_ �Mɢ�G��ԝxH��|�,�~�{T{8��)���H���)�s:=�nܞ���YÄ��"J}�����#�_��-�{��ag�l}�Mz���c��'��$�3H� ��˾�����t/RNl`��j.�	��RzHo�V��TY�ɛ�8s��L|d`�&���#y(��.��Rf� Gֽ_l�m����P)!-��#��9̫.�b@+��st��E>�ggK8y�NPnpK�Bd�a�u�����N��3g�υ�7U�>�v5&�~=GL܏�tڮ_��Z�,�/7�2ҿ�.fU�� *���vH}/ME��X���C)BހۤjaE�� �Y6�&#�yMW��S���S�9>)W�s��r�#�p)	�T�R�����n.�+�����HKg�o?��5 �z��2=0t�i���Is�%��gTb�<���W�p)�j'q�����q�S2X?G�+��9#I���u	�&���6�K!���g���!������Tq�=�Xl2?�dd0l�z8|�a�9�b�~6�fQ\Ŏ��T���7���4�q���n����Q&�Q���'�b�ۓC�i�Nոɲbh�-�L��z�ޱ�U0��q��A�H>������*(ᛠ-[QN��Y��z:��k�%ނ�[��GE�����4��1텘?�8%�-�\��.�d��p5���-2��"L����h�텗���z��5|_K{��g�ev,`�]#� ��%w�f����L=m�(��F�Ȑ��7�V,L/����p��Vt$i���/;kis��;��"f���O�����0���m��
>ݩ��Qr���8�j�+�Ҏ�!*'��)4�=L(Y S��XEq�5mV�tX,�
.�+����*L(�\�͔Gr���ᒔ�&�~�M��j߬��O=����A��wv�d����֊��*/6��bUƪ��+��<ai�FUK��m��x��T��g��s`�B�ް��
;]`���H��ݶ4&��W�(u��Yo�U�Jo��|Q��4*kx,��:Pc��l4���`1�CID-�ӥ�{/s��z �ec��$��^�������~7N��>[I�!F�O��G��n�	w�[����j7�����\JF�Z��Q~���i�����zS�EE�{�F>9�ş�)|޿�_^�����1b�eڻ������Yz	NG�,87���ѝU�0�,Q��!�xGm��5�.5�{f��لɅ<f/b��M��e�L�#�|:����H���mZFb~��̔|��U�\_�U�c�}���xl�h�@?�s�9�w�G�d-yX�n�iim�2�$�z H�Vc( ԁ��Udͩ�K����C�3�i�ݖXK�}8���|�:�Ƀ���)W�̽Dv^�L&g�*VԈw���|�������ց?�ht�گA2�ӯ�t���}Ld�Ƞ�e(��,��\�03�o5x��o��
m�N'`�~8s*9���
��O9�3�%Y r���P�Һ���G��!������j+# �>JC~6-.��D~�(N9�:Y]����q%�.�k��<��t$�a��I;=�,�"�Iz:���62�_/ME�ΠXQ��hse���Ҩ�6X���)���q��*�l.^��:�n/{��:t�l{X�V��~���AX:�;��(�R���b��b*@,������H㕪�5�B��q�����]α�?-euܖ���Zi{ǩZ�P<Ӫ:�<�A�����rܐ���<�&q;��6���ah�$�-�L��.��|xtM�� q��l��~{�h�Ёu����;��%�垑%[�A��y��������,���âMJ�^ّ�]A�Hyn8�U��VJ��V��@{V�!��k�Uw���3)����DA����{�L�#��Cڀ -��SIZa�*�`c���΢��wT~|V#e��M}n?�	�n�=fT���x��&���[c�����{��6`
�K	y-ᅎ[�dh�N���lG�}�l���Tbb�T��9��z�I�S�Q�^����S>W �S5�׹�P
�J�ϷҮk5��jY��f_O�v�4U�\�R�@��D����p^���V��@�N�$m�P]�V�=4��d7r(4�0����B���~.u.�o������qe�_�YU�,�G��-4��u���vӮ��*sT �h��N��<D4���4w`�2�9=�=[[o�yGkޛ=�����lE���)��Y�8���`�Y�ї<=��q�R�e���oo����[��� �u�����5����[P�	�}.۫3a �U^X(���I>���>��J�[w�w��A�)��/'(x'��GV�uP�q��"�t�{+:
��ݟ#N��덟Y��8-��.�xX�쫘`E�́�T}��.2��$y~w���g��_����4]�f����3�ly�"A�B��G�_ZÛ*Ha�������\�;��zό�8��snӱ<��w�ok9�Ϫ�.3ԩf���s6U�0�(n!U};|�}0�'�����?%˗�>�z^�/}���_�~*�I}�'���!)p�L#P��v�Q̫5o��,@F�L�4�kT����wL~����fD�1�կg�n��֟����$譽�G̏���(�!9��4'��o8��h�t[g�_��4���A;���̬7�q��KݔE|{��r�ekf~���w�d�>�Ů�*���Ա?��IynO	��rr\�\��>����p+b�:X���$?�#!�o��'mZK�;6�ݬ��>�	��AAP�3bo�X_@G�-�[Z�#0�	
;�a�<23�}�uֵ����e,�!��mv}ݷT�SM12�t��;�@>s$t��U���W��Q�!J�_N1#`�Іs؄jM �&.?������P��y�$ӴM�T呐�f�bz�XMT'<,�)���spqy�iL�������Z���\��F�Kt�<9I��r���py@>=( �<���C(B�B-f�#�?�O����d=�0SC�Aw��.n|O�/��^��x�_��<��)y�N����߁4�ͷ �e^��K)M���$��>ى[t-O�x�u��\)u3r�(��EG0/w>\Kߦ���E	D�g�{�gl����v�����˞�Y�ϯ�QH���@���;�dN%coߗeB�n=&+��'2OP~����!u�u8��5��h�bO> d�7Dɯb@�I����RrP�\Y �O܏�8��-��)hF �ah�f�Q,4���/� y<�p��4��;�t�=i)�J�&a�c�Iص9X�;>erт�ψ�r�+jdVW;�3��k��̃��c��֓�$}������C5B�ɣX��U�Zc�;n!쭐0l'���pf�4��\�����m)DW��_��ŝF��IVV��\�ޗ�1�V�V6&��+�ʦ��ё����M}�x�ή���s	��Cߧ[?N=z���|ʝ���R�=R��k��Z��'�lj�Wo���B�,2Z�������gAF"z]	O�M|#��bb��Nѡ�w��T���tB�Ne@7���y�y�J����_����%�y�$�A�F���r��J�NY���k��	��y��(�|�޹��05։�.l�-+���d(u3��y�����]�X&��5��R��3	�,+m�.�^��\�(E�$�ᏃiP&�G?�c.GeU^� .���,�oeW�?�XE'[��>�"<�$]��lFu�5!V�����3s��Q�T�3��&w}��XqA�
�5��(���O�p���/D�C޿�{��H@g�U��*ku3U�)�p�{!`�tuE�ཪ�B��7��4epi����֕RO��R67�9� F	D��Ng�_إ�M�w��)�s> ��l�l�lU~�{Ttr�9���O?a>��i4��w޹�����ox{�6�ILH)���Ϝ���N�X0mH��ܵl:Ơ��A�՝��"'�Cv��uJew�	oe{�+8Գͨ�W/ڐ!i4Ee+w
i�lKE,tZ�X3�b.��d~;?�E��+�iՀ�n���г�.c���7���%���DΕ܊�[��� T�bC��ۛst{)�Σ-�ɣ��bVͻv@���=T;]�P3���,F�~���D��zKj@(�(a[*�}枑��4��u�6�ڨ���q��[�[<UU}�W��Uk0.��db_���
�r���.�,Y�V�{�\	N�m�<3�B�٩�uE�f�]u�E�Ձ�m)-��j^��j��rz�2X���f)�徆�J�BS��Y�!ȥ��5��:�evY������o�C�G�~N/` *��K������b鲂|���?}��� ��Ș��0���]L��n�,���ti8ky�����#��-��L��ڂ7�vmq�5�3`%����t�h�QB��bcc��Qe�a!�o`�GT�+�B�����w5J7ܟ�hn�?U�j�!��_n�!*QmG!��M������g���>�v���E�dx^��!<�h�U���e9�sW~8f�g���s����z���wԨ��w�����s�w �P};����J��?��+ ����r"P����B���=v���󗲡Wc�g�{�o�����뜶0�������@O.�����L�^z��'��8�z`*�S�����({x=S� ��n���A�8�<��Q�j���s�'����4,�t��9����B=�f\>�A��jW�����}��l=E�ͅ�J� �BtW�G >�ӆ� 3)��ad,�>�<�����;c�UvDw\P�C֬�v���#��l�jbU����	�֛�H�3��������ʐ|�a�4�]ӨZ"�Sǫ�ܡB������	v�����gbk�f�<�l=�U�����o�B����:`1un� uR�k���&R�	S7�'�D}l(���Z=m����E[��Ө��׶�BO˹�UAj{d�
Q�)��+ӭR�����(۷J�o*m��\y��+����J�$z�c4��s�����q-�V�/15+zI�%{�`�KY�&w��h�!�c��^>F�]iSR���"1ޝ$߂3����۝ԟW�J}n'H���Y�'��4����%���K��FDsT_��v�(�-Zd:U ($���9|S�X�`���u)y3��Ӌ.՛.�ԛ2A��?�T�-�Z�#��1��ݔ���G =a���>��;��jՏ�����B,e+vբ4�r;i�@ �[;�Dqԉ�hZ���y�����\�g����_��E��Y}�ܧLy�A����Ν��	���r�SZM�8i�!�M�+�{ 7W��zH�����dm%}��lO��4��!x��l�(KjpFx&��:��7�>���{���1�v�����tM��l���_�W>�l�Z�+������UE3��+�z^�����e�䳀Z�����'���S5+�c�]DI>�Z�^X&��*;����>*2�D,��#,@�G���b�K�^�3R�jn���+�����Р7�4����[�o\�9�=���7��a�l�eu>�rGu@��8�k���a
f�f�=��:��̗�,�5O�D��sG�22	��;���N̿��Q�I<�q����cS�]��! C�[�&^�f21 ��}��J��Yx���iC���=ĖBRE~�>(B>.S'54��;7�ҹ>�ޡݎLF�=;3Q|��{H�>i��B�{4�	w�X�c���|�/ff�Ӿ��RZ��n�c�_v�����{�;[k�AU����� �Er�}����¾�ݮ�|QvD�{����M&������1�M��� �|��j��Z�JX�ʗ`c�K�H�0�i�ќ�sԌ����W06��&�V���G��`����F���:�'�'���0�EA�*��ƕRqv�%��DUT0#�-H����/pE:��E �GV
X���5���O��t��ֿ%�����U���=�K/8xz���5Ptю]�;�r���`T�� A��-���ޡ�W�C� �U��k&�'�p�Б���(��u��q/�ˌ�+�Bژ	��Z����gx�4����:�+�`*�j1Z�VXw8u#5�n��ϾO��
��ϸ���?^z��S�w���;N�=t�O�rZ�)����]��*��bd\:ܻV���n(4���c�Nh�Խ� �$�o�yj⚑���K�yW�y���N܃Iaz^;�lݟ*W�4W׸?<�0j:�5�߶�n?��5��٩B���T��aQv�׀��tK�H
(����H3t� 9 H�t#!ݝC(!9t���Q��w��0�u�>�����k����Xt��z\j����b�_t"6����^w��>5ol���t[_%3�1�u6�B�P���А�����x�g�y��%��^��<��{P{��T��C�v˱�V��Q}��q>���\������F*� ��� }E$�#^� I]�D;�:
qǨ�'/�&�����^s�жZ�J��.-k��
�D=���_� �{���:G��c�����/��Rw(3zg��OQ�c�kl��}Đu�������ץ:�`�#�W�!}��.�hHD_�6\Q������ƨU���i<
oK�rkk6:���N�'>�K�z(�)d¹��G������ss��[l755;�x翡���p����5 `{k��x�ި0�gz"d����S�D�5N�9Ws�A����g=�D��I ~e;H�C�y�@ȵq��Ϯ�f�Tx��ZR�Q�{�:/�;(��U8x&i��&�`�`�u�Xஸ?Y��bLjP���V���_iN3��r�>/����k��~CÜ+l�U0�y��x����n��E�y��&�[G^E�Ƙ����ۘ�0�!D��m�^����{c)������2E΋/36I�)Қ�O���3x��+0H�B>��|��oH5�Lv�'�Y�G�-��w���#:&�5�ˈ����Ɩ�C%�[u8��B~�[��xW����AF�f�H��%t�(�@�amd�p�z��Q�p��Nm����������mj��˦4¥S�B��:�n�������%����$���U՟. a_,33��:q�G����c���ꗘ(�x�_9j�F���Z��+5R�U5���� �@U���6��k�cUr#�,1v�fEd�]�RM��Mxv�BZB�]�_�o��	u(�����J��>G����n|.���_�+
F4\�exa2�)��
��M����~���ֈ}�fϞ�
����%r���~��e��?=�Wn��%yմ���=�^b�uF�-��c�pѷ���#;j�!j-��t�m���%a�D,�:�Vv���T��#��b�.y,�0����qu��{��(�?EУ��4R��:��������ߪ���@���0:Wvl��yf�~����i�")�� h�}�b��3�M���
�=(h�:XV���F�����$�Z�*6�,��`/V՟d�
�+0�p.*�N�Iu�8A�]�ԿK}�IU���Q.:��}��������{8�|���nѦ8$��X~���E�������u�/[C�<�5��m�5��]�к�����
�꩒@o���`V!��0}�!��������u�Iª�T�j�* F��,��%�dHEɛaEH���U>z	�!.ׁ��8}v�q�s�:���\��+��hi�b�$�KvR��52w#	�RQ��>9���Qy����%��=J�i���������LB5��¥xԝ�iJ[�MC�
vo�S����|:��

b���鮜�@�f����G/��j.�����5�P��=����I����e���^���i�����@��d�,��D�5��8��H/�C�c�K+d�"4�y,qʉeA�·���](�&��X2O��I`B��8Q)�܏��O����U�:'c8���	��L�||>�[����p��Nw��S�.�BuH��쑲���c�:?�=� *j�����$��\��O �d,/!F���]<e���C{�KZ�eCܸ��x
�C�g�{ e��?����Q�"��Х]Có��w.�J*���/X�{����H���}��!�o��gH�<�Ӗ@zܧ�׀��dn�^�ϝl���4��@�&"��� y�X��`)79ͥ�띶Kf�a���Z��L@���wU�Q�G|���N�u��v�L��lD�Λ�w0o�y���:u�U瑙���R|㓼B�C��Y�h���<^j��I��:-y��� s3�U])/����*˽��.����h��@}�k�sjs}�E�/w�P���7�Cx���U�Z�h֩�r�8P�_S���{Z��F�#�R��^��b6 �F���*�?��M�DV��1O/-N`?�2	(��s���7P�ϛ� ��n�Y��<��j���=�/���#���|(N�����%yD���I]��#���ભTδA
��Xuh�Q��;��
��?6v��\ܙ�G�Ǹ �E%qDݛ��6�KI!��RO�~�o66G��+-�j�BSˊ�s�6g��]^�>�֡�XH�:��U��G������'|�"ȷ�[��Y��-�����7Xf�\0k�[�m�0��c�$���=���O��L�<�K�e��9՚'����6��k� ��~
�I;C��ڥ����^��unHT����9�fJW$����C����k�Ul�Ȯ=�����獝Ǻ��Ĝ�R���������xa�m|+��>��2�l>�6�X���V�cg��_���k��e�R�X}��]}?��J>��Ǐ���}�EkJ?)�Ia:'��c���I`�2����z�R�B����}d�c�<�D�"���_q�<����~˓�"���͈ܳ���<�bQ����
�>Tuw8�w���v>(�:.:�~m��w��|�jZ��Ag���t�`�-���w�75��.@Ve[�")����X�ݱ��$��3�-�gB����)���jEy�D�G�v����W"4-�[)��b������vI��)�a|/�jj�]�#�F�/�nM߷�<�(�ț�qH��:�ѐ����0��.֨jR�UZn�g0#�q֠�O�����1�0@�o��J�+�\{��G�QS��"O`bz&6��+u� ��s���Z�L�KHR/ Gg����K4�an�����O3oq���202;�</�A�ǣl^�<�;ꖺ򃧇N,*�W��O�����`��iޢw�y	,��(���3�i���>~�G���
C�2�������H��e�Az�K�.}Cv��x¥c/�˨	8çb���]@��FI�92�.s�C~a�V$R��bf�5;��K&NSZ �ſ{�M,�\$u���*������m����fՠ#�4�|^jm������m���ׂnK��`B%�VV?D�ٳ�ҩ����=���֝|���'�u� ��o��g��N�Lx�(��*铍��f�;�Z7�U��0$�7L�^O ��f�&)�e�;x� ���5t��wI�d����ㆼ b�_h����Ej�4�˪��� <H��OGLn��_�p�闁��(�0�4���"ϲ�t��5�#lM>�zf��E̖6�$/���;�����kt��
|��C�!���������y�Ă-H����qıҚjQ�g7���cA�p	D2De1�|c�R�L�(��W�~�~�\�� v9I��(��w;�R��[OFTնk	9�.1<5��`�,r:�}�MA5߻s�>̘��B�"aߏ�)��P�Rտ��)3��?B��y�	z�{��%��`"�I���jg"�JCy�G%�dB�R�Ƚѐ^���j�Ma)�2�щ��$���Djm�ѭ�P��(ʺ�d6��%_�r,-��y���Gi3�q��=Â��kF|I@w;CO졏�b+��D>f�)L�� 8���#%s��'��oX}\�@�ET�'�?����>��ἊSKQs�K���}9�ɘЄh*���]E
՘
9ەt˸�I4�s�GZ%x�-�[�x�y�e���4H\H�o�~�#>� �&l.��˧8�}D��Qޖ���my�ǥ�J�`[��{	��J�Ӎ��0�ˎȤM��Ӂ��b(r�k!y����z6
՞�Tܺ�������/U-�1�]I�#>�=4ʭՙ U|.������@>I՘�E��°Gl������}�e���5-5���@ԥ8�e�w�m
���D�o5��G~S�qzފj��^��L#����}�bǌJ��4��$?�ټ叾Q�x��4�^�}ފ(I��oTE�~ƺ\A*��]�=���3�|e[�yM/��Z15T�N.pW�Ą���G�l���y������Y<\�X����f�T���&D(��s��ǃ�f��|�Je/=N��~#S��PDȎ��8�?<q"���%H���1������z*I�.�/eP�;�MY����#�A�q�yW�:}���M�ճҢ�����®��(�fiy�\JiE@�j��ogw���WG�G �\�K��;I|p?y� k��դ�f\aKރ�4	������_<з����?M����6���/xN���z�n��wD�f�@�h0-2_�C�w"~�&��Om&*�h�N�ECa_>��N����_,�6�svw��/��
 �︨���/}�(�-�P�#ܤ/�D�O���j��,�J[�>Y�X�-�D����*xT�@:�I����f�SU��:I��>{�vI���s;qx�W���b����-b%Y��2���^}�{Z����NC^�⋢�c~���|Ul4�+�[�x�3y�,�?�w�~��q͢i��g02YW��R�W�u�U�ݭ��w���EӶ�y���o��h�ˏ>�Gj{����pk�ƞ\0!sI�C��a��o��"B�`B�8tĥ�p���9����׹Q�����zKx���
o�WSQ���7�Ɔ�5�!g,�3F��!��2��͕�A�Ջ��F^����e�V��^P�L��n��F��
]�Zx.3bza		�w0����.��t���O�.�E��	���)ٓ�pm{r7�3Qe/2c4ur]�Y.R��[䄲��������'�ϱ_�_���/���a�=[gX�}�/�(UӺg����84B��� �r����0?�d`�P�Ӝ��
��2fq��Q��/���\w$!3t��@�<�o�[wXZ��i%<��%.e�<U�ZK�W}�ϲ�:whO���Na�H}'�2�.nx���y��g�BE��hi����/��h��@���^��(C���s��4wkG6�h�i.�h$3�ES��=���Z��-��G�iIN�N�Kzf�����s|w��������/&y��R�G���Q����wK�X��g����H9#��{�xv{K�x)�����̢��z���jH�C!�a��w<��Ҕ�Ul2�ژT�b��C����!{8]�:���CfK���R����8$lx�\䴺.���*S�c�v3ٵ#9�)m~�.�㑒�����¾��˅������y��/�������u�M�{��(j��}ͱ�BR�{h�N3�DQH,����=)�����i�gql�fa�N4��T>���q9�=刵$��Pb!���gT*�H�y9O�����w��F�|�������h�ږ����ުӊ��@��nf<��d��8�]T�G3���Ҙ*���1R�ti�����5�P{�J��{��L���gd%�bg<��Ə@z��Vov�����6�5���	�wG�c�\�/��H�ܐ�V-��k9���ʈ弓P%Z�k�*'C
���0��To�!|�)5��z��ċ�
8?��F�7�ahu�o�a��s|��������"J�p���{�iRKLQ��Q0�>Sm�yN��Bރ�%��j'=P�޶�7�f��b:�uq��E�;�|FT������wcJA�?��z���|1��	](�Jl�rx)��N�.�?��j})��b�}�l��f������'�N<%r�s�z�'Y���Z�.:� ��P���)x� ,o`��9H#Z�F`׻"���r�y� ��kr��E�D���O�g,�Dc4IYF꺜��~B�{�hθ"��m-ݻJ@U�'�!ң�_=��@f��e4�Z�R�¾�e	�}N�	����R>�0��}�N�k�eI�u�9}������_�G����u�U�o�æ3ō]�$��N����A��q$�$�
�R)�ENj<L*<�6�Id��fVM>E�#�������w6I��O�͉}�b�J�ɦv�
�	�dx'���3�׿a��u��n���6�z��;̙�ϖ�5���B�C�+]�:wW�~����L:�c�ż2�qe`>�`��������y!?���gv��(��P��oO�>[���P���y���Am�$׍�ۙi����V��h�j,f�B�ё}��K��xC �eǆ���A�����n^�:��> �F��x���n��ŕ��H���ۂ�q�oʋ��sQ��c�z�����wu��-[��g�ªT:0������[�17)o�ͦ�9=Hȑ�u��g���\H���������{}R���Eۻ�l�)��Қd�$�9�Ж�n�>i;�W�<�������	�
m�m���	���n@��Ė��9UIy���%���(Ր�g��
���n��/�f#JJ�L��i�����G}����b�4K�WWW_��o��X�٭���A�Ȣ���Բ�}C���ܿ�r���o;�� h��Ѹ�w)��~��t�m�s��y!I���I�d�=w�4-
l)��� {n�c��)����}�1��o���cki���2��+���L�$w*���M8�}���@c@��v���Oh���:�ռ�?ɄC�M�5mp����bJZ��c�q7Тc��;�wUOV�1'� ��ήm�~�@�1UA����[�Ǒg
nZ��3%�|SxD�>E�Y%�{^��+
9�fR��0!�ª���}xxx~�ױ^��~nj�oIff��Ű.62�'�ǿ�����������^�����˵�|�-W�"�}�9�F�6NZ	�~�۬;p��MF���BAy�Pc}N^ڊ=�^s�u,)��iXL��1�?e�
�m.Jr�������d�9֞R�L�]�قFBK.�iF\tb��9�<�u���,�Qñ3�ɦ�i�cI��"-Ɵ���~���]x�@BA��F����U8Sȋ�WR��7P=M��{��;���[E/ɢ��x/�\��Sҗ5|�����T|�ܽל�fTZ⻓1�;�O�V�:��P	ucb')@hW�ש�����CzMD9I��w�[���#KEBT�»�C@��>NnFa�%�Jx�A���E��ѷ�zzQ���|�ͥ�)�8�5$�`A�`�D-�\2��)!?����m��K�]e>$EGo�r��$���Ml��"��J-��Ը7pDVʴM�ӛG��!����J�0�s��AN5���bCR�����Ql"~��KfRm&#s�.�\�ȃؾNb��ι��-�����ٓ�q�w��4��~e찺��"�=#�b�f�a\���3-��\��}6������/(+�TE�b��Dn�.������c�:[xLZZ���Ni�g6��/_����M�.������h%�����]q�����R��~�j��o��灔���$�8�!�i�9�i�]V_��~��"|�� ��:D�aeqYz��,�G��jZ:����]��q���K��>��Qag�� v��tㄟم.M�3�|$S0ImR;�xl��o�б�ow|��z<�7iU�����a��Z��g/�˵B����NM�ѓ���&E
W�<�ŉ����޳,ˊ����[��|g�A����k�����5.�dwc�Wg%껲�F�W��� �d���Wsa~0��� ��Y�lW�H�����o��*k.��(-\C�0���5��Ԯbo����K�޽�!n������+!��Q���5����2��-��W�@Z��i$����,�X�R&Gb�w��tQ�����r���l����b$~�e�c��VΝ}9%�����L6*Y޲RD6�� �r\�Ԍ�klޝ�����3��92�7[���6��H�4��o�#($���~�����F�vYYYQ�U�������_=�v�'"�-�}]� }vi�Ŕ�>ʹ�ǡ�'������)7b�fb���7�r�tఎ�M�p�^�D�i�}�:J2�r��'Z�{6�7I�&Uo�8��B(?7�X�0's�cN3'�U5"t̫h��~��AS�	ݷ����8��F�J�[�"�[裤���~������~��v�W�G�c9��A&��+�L����v���n(���u�[��*�x�Nf�$�?��E�ҺAKk�(�0)ro�V3gk�����F��zo8�=I6�L�wM*E��f}��^���j��[�]&w!@��nC��r~��|��[(���*�Bn�[���Җߧ��+=,�F�ܞצlI��XǰChZD˃	����23p#G��\���e�xp"�m�jx�j��M����K*�υ<Ag^ї��4�"��i�@���e�;��Y���:��w4��r����%D+���=.i���Ì���u�̎C��X���:���@n�Rh$�1����;�Z��w�gB�K��փ��%�:b!�%	˼�>9����A� x�>x?��Y�]{�����O�R��ly�
RH��c�!Z�$���SC��*\�_���q/�lD%#�O�k%�O!R�\ ��sF�2�֛>@ɠ_������='�0�/V�E��%�֑�������_��=��FQi����o��YP� ��?����12toc�zq��k��iV��薬ے��fz�I�y�t��O�=�����NG<��[e]���Y�W�|[�E�N/<�n�)qW'8�_��1����;sBP;b].O��u�JR[��*;���m��صDX(|�h�8�rjl�}
<�!��_d�w�ŷ9��_�ߨ����W�>�گ\�� d���T��k�O5zNj�-a�΃�N�Tŷ@$t�-��H;����l�zC^��C���!ma��lnԚYl�!�|)��R���Ξ~k�}`yR���+A�d�G�֟����	;�	��M���JBԜUw�#v�Z�2B�/�z�[vG�e�[�K*��;��q����O5k�-�{�fid����ʴ��hДgF�,$�S���mS��h��E�8ʤ��i����f�?�?�,]�V�߲`D~,�����p��w���n�74�I�����?�[���g)�tZ"�M<g>-͗���*s,X�s $�k�������m���_P-��o�m�GW���i��@���A��qA���!��.��~B�
��y�N�e������I"$�S�="�
u�!�O{���M�ȩj{��4��f��sJ5�wg�HG~m$�յ$̬�T��&��c���Z/8���lq��e%9:�h���[�M�d����O������|Ugx�<`u�)�O�>��y~���m?��4�����l�R���JĴ�~����]�J"��X�l�J�nx�m��/ 8�7<(|���u�;m�q�nQ�)��vX�ܫF.|<�)F�<K߾���g���
b]�-JV7���x������D��W^v?��<5&2�Oc���E���;!����u�>���i���p�D��V��Lϙ�Z?&��|h/�Ճ�Vf'ڰ��S~%&θ�
ёIΓ��Ť���+N��]�B�r��|%��Zi���J�@�j�ҩ�qkn��ZL%Y����N��`���i3���)�J�^��@����f�Ebv4��fL�@e���8ٛ�u"���Y�[Y�ݦг�R�/�_�C�Q�'�ݖ�����@t��Ϝ���n�j�g,X� �_	���6�j%GҾ�Ļ��J�v�s��~d�de�6<�Cr��=f��c#i������wY��tf��~�.��ɀ��UNd��m�H�`�y�|�7����t�o�Do<�H�����^OW���'��^j|ɶ��W4���ATu$�2�.��;U��y��,Ya�-���1?�ˋ[	�����&��Fz�o�0Ku���y����m��J������;�(Y��T��~�v�q�%;o��w��Nt��G��?�HD�>�wK�i��@�^dw�.URQ�y�eb������HY�n!>q{cՍ��\T{9�]jS�R�G�9U[P��\Zz��]?F,ۏ�GX�]���٣��g��Oخ�̎|�:��Z2��b�e�on=�\�S�/�N,��u̕��巻�]���a��gI8�"�6ꄮ�j������<�\��Gk\��B���fq�U㆚>�٥/.�_����iХP�pT�&��-�,8Y�c�!E�����Rf��= �;����qp��TO�
Sݦ#!9��і(�M���^nDtBfz(��Y�e;�2bW�N>�s�����y�0��ة�w�:@�y�:����9ʮ!�p�]rM`4�	�-Tۆ׽����(6�U5c�_S����B��/si���>��r��o���(��$M��8M�h�v���mVoa-����(>��XA7�	�6D8i��W �W{�e����v8�|ǿ��<�R���كL$n�i��nh<.�:N�R��Tb{�eM&:�c~�c�Y���׷�4aS�ꅄ��¥_E���Fş���#ABz�1���&E���3Ya� �i�A���\N�MgF�m��R]l���[�R3l?R.�1���r; �b}��oI�yFC���?����{3 ��\[Y���Nw7e�W�� 
[�۠�<��xi�w������j��ۦRB���	�q�̬n�
�����%r�p�ћ�Y��5�|Hd?���
�vjn'�	�i,i�^��ỉ��Z89�4z>�[�>Y�H��p#!�Gc��158>-ĵ+�0��-CFB��rNzL��|�k9)aJTL��(|����a�h4ۡL��x�r&�|%�溹T�">����Ƨ�RSQ��TTZ��~�8@�,h��F�l�jT.�		�ӹ�K�_�l�@�a��{����WCB�$�~J�V3�KX� tb�g���rNԡㅸ݊�9^��bx
v�]�=�ee3�@��٬uR�j��\�f̫��� xugy�<�!���_��� �h}#Ѧ/P0'�<xt�)x�I��V�-^F_������4��aCB���P9;��,��0?_n/ٽFmߐL.�?��5�r��;����r�7��f�B�Z\������䪢JIr��jlO0'm=��*8Yq�VW�/�>���J�q�t�w0<(�YodV��̻:�}�*ў$��[�:�YX��ܐ��/��t/*��&��Lx9����zM�|4�dN���h���B��ĥ�oa�#�Y����k�Ǖ���'��|N.O.���]�KR;y��|{5l�z?�x�Z�����n������$U��&�iq!���3v-#[	t��tu���C�D&2�Ճ�<g�.#�y1�i���I��L8�I�־&m�����ݜC�DN���*�z�X���s���\�8r��x�B��� �`���|��ȵ����r�������:��z��!��Z;P�c�;�q�~(Mg�c��ZFᷟc�kh���J�<�'HH9Y���Q8&�-WkPcXee8�W`�=Ԏbj�n㷙�T'�j)IXH0w�
Y����i��� d~�$�j��6�:�KW �y�#i�Ey�&��#�방��&Zm-��\M��������^%�o�9�����[�57������$��^�La�)��J��;��EJ����ȊH�K��~H�f���b�(�۶�*�����v���ULdF"����1�Q0m#�2T�"�\���@ʢ����x=�t��v�FF��Á;���[��a����f���K)�C��1�?��	Ve�n�Y������|�q6A8�d��S?�)��d�5�xXŧ�:�S��ȫ�#�4�5�d��)_����)K��xC.�$�r�3��S���q�*E�j:�/ZJ5�.1uA���W�;2�`�) ~��Z�p8��'�U%�����Kf[],�w�n�s�]ƛ%�a+ku>};e������@���)�|'&E�� V��h��w�;x5��k-|�V�݅w�"�
�M�R��b���w�:��Y:�/��?Ўe��&CS�����2f�����Ζ��i>�Tk�?�_�����M.�}8��y��c#6_�P��}8�]�=� fѐ�%����ګ�zgw.6�
�� ׍-xc�jղ�T��W�n�(�LY��;C��ܽ��G��"�R`�b�^�ՂKk'�ԭ�[�]e�:�&��S���v���������׮�L�Ԟ���QK��N����+��*;�T7���MB���mm�2Pi��"$�K���Y4�hm(Ť6��nlY#|�Eft�����a����Z���H2	��Ԭ<��V�E���Cʷ�
��[���oeׯC
��*U�b�X�(�f���w
%<ǀ�#%0��'��gZ�����'�)�`^�<TSW�b��yr��&m�&�.����՛����S_���R���"��y�ȼ��⺾�G�9M���b�i�����O�翩Q}N2M̆�� �: ���&��uem�A�r�.��A�!�1��"��`�T]g��#�܁�	���Ce� ���i��$�� ��x�yg�W��ũ޲��e_aI[y���b���K���[�xgl+��n�qV�т�kx�ʺ��I�:s�еC�!��x
�4�K��x_�n�]�6�VU��k�a2o�:_�v� ̽ˤԛ1ki�WϢ�K4 ��Eؽw�E�>c�J��4)��p���c���s���k5e���E8$!��J�m�bX�kIZ�_�0={VWg��d���^�ݨ��%'��K7N�MG�&c�:�@_����<��E�'G������-�[��}�ɩZ����A����/�0�T�Py�f9��E���c��Kp͂{��+����{��z�� �p�[�uf���]�ЌQX��-k�K�OK�
�������I�q��mf����=tsZ�ҝR����m����Z1
 0���ȨPQU$$4��� ��A�&F���H��!���n��C���9<��3[W�+��-+`飯��X6CT�F���h�>|v�=)���x�;�C�������(��Z���4��c�3n������|l�!�;��lu�&��b[�e�5��;��$��tq��Yɫ�o���Д�o�5wc��	|�:�A��� �F�n�,�P�����w5w�T5�濺K��T���<��S�O���Jꠘ~>�:�էo���}5���ֽ��k;h�t�����G�r��uʴ������ez�������f��4��	���u4���1��)#��\�^:���t-���ܬAO	L38@���m�*����{y}�����ǆ�Ӑ�!�*�E�M)��A�(�����k��� �s�C�w����&�|S�$H��M�x韑�f�4��gi����p5v��,.~aޘ>�av���Csel���[�u�2��<� Q��<��b����ȕ��%g�=\IFW��w8`) h�ӍD��#���YP7�^�2�z�SY�Y5���5͖~t��TH�p���oI��>�K��m�������ԧF�(GT�Y��;����.;Ti�y�֗�N5�k~�גuQs�m�݊�=��m�Ե�|���<���gх7k�|s�eq8D���'�k�B:eT��z�1��KT�<��Q�����?S���ki�
k��ReE�@˰�շ[�W-��B����Z}�ε�p�G��1r��l@�$[����M�k�.&w%!9I���kP �ӿSjθ�g�����M��_�Ez8%��L�� �x�����LM: �{��E!UI�2�&B@Rl�%�"p(=y���ܻ|A��kI�i�g߸h�F��ǺN36m�����F�p����(��qX&��#+���\Uq�a�Qw�f��Cm�1/��#p*���{q�(��p�����dC�c��V�xW��6h%��!�+x��~9}�s�e7�2��d4R�vPF�tq��]|Lr���g;�=�6�ރ�Vy�-�G}���WDVTҗ�x~�[��f�l4_��q�[�]���/^�?]3��D�K�,�xM��椆��y���t^�����{�Q�we_�1�@�ql���2Z��>�<r��L��Z�����N��8��r7�4�Hp8�qy�^���7��1��^�����V�����G$����Ԯ�bE�Fl���.����)�I����T-fnM�xx���_ 舭�JL�]���.H�:`�	�A�IH {�!���}-[]+}��	c�S�����v%B�� f�5c
��ܛ�(d���l��%��4��;������an}-�3�mp3�0�J���x������!v`�3 ��/?��e�������?��9�!�޿gh���}���||��h�<���?%��D�PK   |��X�ĩ�xa  na  /   images/c9c0af01-d4ea-463a-b9af-0ddeafc58269.png C@���PNG

   IHDR   d   �   �oƬ   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  `�IDATx��}|�����ӝz�\d�Wl�ml��!����蝄�nB=		=�б��ٸ��-ےe���m���=�I�fɆ�?�gI{[޾yӾoތ�PSU?���ǆC��_�;��OHQ�^��#����k�G�X;�����V��hQ�c;�=X��� ��c�v��?�����;1^��d������(?eohd��A.��%�9�?;� Mރ�!xI;̫V��VZZ:pԨQѼ�<Scc�����+-�����LxF��9���jZZ~W�������s�T�`��T�_�����S<���P]]��~�-��۝b�X�Vr8�����}��%���5K�a�����N�M[����4�����t���oG��f�q��l6[J��������w/�X��frgܞn����٤�-��C$�m�y�~�8�q�ܠ�}�O�(m���8����:��
�e� ���s��Ü5�|�j�?|����ZŅ�s�y���͵L(�h4*���܃�ᣋ���ñP������{�#��7�s�u�!������_Uͳ��!���4l��XC]�SO:i��{��nQ#�ǭ�Ǒ����w��HE��]I��똔�I;��ъrRxPc�dr�S�l���G��2���(
�\��Dh۶mT^^N�~�)͜9�\.���4�����Ӛ5kh�ԩ]1hР����.AZ�������Cٵ�@�����G�����}�q����7�@*�WQ�vf��m� �	S(�?Qx�f�HǗ�C\�\H��A���y��`��4׭�8������gC>&> ��͛i����EpDCC͞=�����p~BL"L8&���ٺ���R�����Ea4"�0�/!Sv�^/O��kn&�n�*aDDZǟJ�ߒ����3Y���z>���a6���59�9���v�����t�;(�
b<
��ʔ���DL���?�G�'�|����d0��p�^x��̙C�{�<�Ν;iذa	g*�_�/�h�/?��ןj�aj�m1,Ń(�;�>�(�*�[�l'��~������jӅf��Ԡ��<c������~d�%�8� ��ҍ�][��Hq�;W7�M�YZ�~�_�	��N��¯����۷S����EE':8N<�\�RG�29�yQ|������%9�=���<��a�q˽d�<�n�Vƭ#��ߙdP�?�Y�g �0�̱d�5Yh`}�T�6�H�\:dM��R�DW�j���dee��2�А!C���9;c�Z�n]�q�$|�$�Rv�}b�"�|y�����I�>mH���O������~�5�L^��x��V���T%u�kv�<& �`��Q|233i����k�.���tҭ��J�����݆g������$\a�H4��k�A$٧K��"
�ZB�_\��Fs�yy^{�bU�:]B���^wsH4I��a��I~�t*D��S)���H�y�M<BײE�B��ޏj���l�FX�F��s�)*��n�����pG�� �F�I˖-��!��I4�(P��/��ig�x�� �_^J�	��u�!-�ᾭD�)#�,��)�w�f t�Zl9���l�)�f:��)�<C��-�Mb�ׯ��w_Q桹�y��0���q�����iI�`�@�HO�ie=�v�yV7d�ƉLg}5���%�i��Xd���:f|�pӓ��8d��(Y��暮8�2z�>�>�5���d�Ÿ�ފ�W����%a�[���� ry<5�{3Ew�9ݚ(<ȡ47�<�TR1C�YުJ����X�-o|��/�Y1iy�4W���k�PFَ����XL���&�NQEM��G��$5 �����V�E�y_u�G�"KD���R�1t8.��x���]�+����G�#snEvnc.I��|�I�*����9H�Y��Z!�:҇�����q�U{)��.8�v�6Wd\sEJ�Qp���i����.?���EU�=;)���O��Vi^5��|��K��I�5���֍;��&��g
QҺJO�a4�쒒0��S����Do�Ĳ^�;�1�R�_���tw:�<�Oj��&�}�;���V�%�x�_u�X���cRYx��?%�Y�y�	M&�\V���K!��ځ��Y����kbH���VVo��P�&�.�I�R7E�蝮G;6 �K����X����CR���*������3￞M��X��|.�}��;o�n��|�Y�M��������+�7L��)8fL�y�� �����'8�>a�>|�Xp t"��an����b^�(u3;r�.z��X�D�vQ�?!�1�x�K3O�*"�b�f�|����+`�ܰ+NR�X:�k�&&�\0Jq�"D������X��P���mC�Lj�׹ߔd�w��[�)���:D-8�ȒN�Z�>�	O��1�~t.U_t�EU4q �$�y���	g��_{�b8�h��a������5E����3�>Ņ!��*�Rc^�(�̺*,�$�?�,܃�b������4q�ZD����2e�-~��j@aV(��>��V���TX^I�MM!�O3���-�����������鐅��Oپ67�1@�[,����r��B�R��{5��G!�6;D����(�1
{���\�����z�!�ȱd�q,�C�[��4�=|�4Z��	2�Մ�+[ D#Vm�!k�%G�@D5�eӒ�0������6ԏ���d�i�Shڧ�)����Sx0asB	-������Q������W:���r! "��ҵX��x�TQټw��r�|��YbP|=����/��'\5�x�K7Ӳc���<���}��n>��I=�9%m��q�A*]�5i�뎡B�cO�i���L�����~Vu�t�)L�W�vk�&>���k�|��h�Sx�Rr��(5�z�̐6D�\ugl/Њ����Qp��4H� ����X��X��g��Si+�p�p�'���'�{o�ZQN�G����^�������wʿ>�y��|��#�hW9���N��J~f���\C�<�{w��%�z�qC��ɺ��d����a�;J�����M���C9O�L���QRR�29��b|�����1(_,"aU(-�[{�@���zA{��o�7�ob�i~�j@��=�,^z����w�{�H����E��x~΢�H�3��i΍���L����R˺�x�8�X����ȡp�ƾ��� ��iT����j�(+,pt�,s�n#SV6��6�1�ؾ
�ٕ�ʌU������<p[�n�ݻvѼﾣ�{,�c�&�1�N���+V��U��c��t6�G�)���ϗ~+�!7�j��}��)'��d[�����yL1�<�8���-�q��<���|���v&=҂>X�V�1�	&�p�y���E�l�k4u�\0T&��5��^b����q;_;Ơ�`��?��h�B�5�Ӗ����Qf�3�ƃ�}G)���+d�����^�E'��F�j�]�'ӡ��SQa����b���\�����%�HXL��5��� Y$ˠa�oEW,!�i3D�XǸZ�a�.�'s?sI�.�B�'6l�f/e�5�G1������ٿ�n�o�@�f��E�U�@�&ŀ��@?�οX`����)��N~ha뜇��2zxv���_{�u�}�@�Cy�z�(���)�u��]�5��\g6�l:�[K^�yi�TlRiBS5}��5�;_��G6�W�h�%Bc�3�/� gj̠���/���%%d��>�!�Yoe%�Q͔�*ں1g�j�%.+���ɚ�My{*e<y�͓�ݦ��w�OX�;��3f�ʍɝ�FR���YY���l�Ŭ#�@�� ͑ȧ������X:7���M!�`�8�M��&�����q�]�����(p�*���V�������x`��I�WF�e�*;0�?�][�6�E�n��Q�:- W�iM��Jg��6U�U+.ؘ���a��rr)�JQ_RW��~a����TW�zaIX�VTF����?!ӐaT�f)�+���x�}���`�Lc��?h�f��$�N�}v�q�k�?|,�l�l�;_��/ba13j�귣<�A�E�b�aג�S���6F��/�p߭dz�~�-�c�G��Qf�ڎEMq��e�Tߵ�~�j����3e]Fc�E�	������>���Yw� O��=B��K��D���RZq�Dj�J7�b�)�7t'&���;i������eІ�SUG��ScN�t�l��ݔ]U��Sq�{��NVR�[������l�2�Kr2����v�`sT��hb����t!|l�"aa�9�=�B��Qx�Z��WC3f͕��=�4�����>�����!�$��ffm��n|�3P�51���7���n��4�9)Y[��My^T�O�q�S�u�f`W��97_|��*U"�o��zX����G������=�?@#VnbU�-�t�=$��� %���&jig��]*�x�a��Y`�����#�t�ƌ�G"�b�
�,�YΆ%Y�`݂�)�E7y��l�/��i��	Q�Y�����Yh�r2İ8��d�0�� ��A{��Iʎ���=���H���k5֗�?� �"���BnM|�5�A}X���kɲr1h�AX�?+��y�e�XY^.���a&s *�ϱ���4b��Ɗ;��P�۵g�{��%��JiJ�����6ho�n��Ԑ�%�2Y���{�3�@���k��Rz����i����J]N�mٺ����<�rʛ:�|��+I(x�⬫�pG���W��cH��&������"�f= ����#S������N���B�U�x��Rr�W��
���J*����5}�	��4��	���7Ɗ'��L;�r���ތ�F�`5�WTu�r�H1��r\.*�̤��f�()|Uߛ���N,����gb��k�'�R$D�ywf�$@ ,�bXeeeǏ�g�-*";_��x[(���ส�2psiZ=m<�+.J����W�k��G{s3i��S)�tp	{}<f�2�9[�nڧ�Q6~'8����::}!���J�=ӏ�̙O��Ĵ�ef�����jz�vW7����8��*θu������xa<�9ܔ�GYz�	R@����x���{i�1���_��n��Y�wX�a�c�bDI��m�0J(jG��X���淕hLm���1_�2�$c�a�i��ZzɝQC�f5�l�<P\�T��)��`{ �L-;)OE,Ժ����� ����/���� ^J"`,]��j E�e�ыx��+ϧ�G�%Ǩq��aw�<����^��i���E��/���6:R�_pL�P1�;�3����4 �||�+�!o��\�^�-#F�)3�����g(��
2��e���{s'/�ba��@0(�:5���}&hMf�>�P/k�x �w(�0+�3�&S����= j�E�
�8�ڻ�7A�+-� 8��c������(+��%}��Kvo5�Di;�,]V�#�˘ �n���O>ok�����o��虱X�-�^�N�4w�����p�P�B|���^-�(�מ�؇oR&�S�zMQ"���`�.����g/�lV��������c��c`�`J#��5��BU4����v�k�>���[�Ą��z��am���X)D0�qa�cT��Hٶ�����}= ��!��w��k+S0-�@{���{X�!q �[�x2�@{��S���d�w0_<�lh1{�^jWI%�G���-�O�ٿ�t���AZD6��O�'w`ᬏ���\��~�__ R������Q��O?>�-C��컷K8�kL,ˮm�nYON�#�i�-,���	�S,���/ܵ�B�֒܄�C=z$�a-���E��/"�K���d8�@{�@��=A�d���%	��|�N�7k09fڂA�;���DX�RL��@s��V��a��.�4���ŕG���C�~2���"s�df;=��KQ6}�6+����;��a��,������kv;DƱ���i?>�p(�~A��[�m����$�|Lm�.��v���s�4z���A��>+�
�a0{��s�I3�1q�;�g4l���3����`�5�a���KD:N�1��Ρ��}T����XCᷚ�3fA���T�� �!�PD�ē�^���T�f���3�c�9�#t��q+��C�la	k�N��4Q�Z<�dYA��FR�ˊ�Ov\@���Հa��A+e�ב��{��j^��7,/�P;��WYX��i'�N���O�dE��]�E�{��fn��b�N:�TJ�8��K���k����~,���J�2d�,TEY\�[C{F���3�]�Y�����ߑ<���{/�T*~^�ժ��f�Y��6L}����bmo�"zd��4`{Y���"30C�]M��J�e,�G���cy�+MvSur�(��i�y�q$}�D�&���md~�k��=�soH�7���u������dXyJ�y�\;+�lW����f�z���ࢹd�q<���"�g��o�Ҋ#'��2���O�`;z����E�$���T�����QB�v
�h��]����������(�a�ch��23anR�ih x"���5c�ƗLU��}~��
z�^����2�����*	���|+W����i(������y�Fg�� a��~u�@�Pd�z6��WӌY��x".+��w�z�Ǔ�hg�(�N�^;~u�SU�8��@�F{u�����5�D�UW��_D��6����-40�&a����4i�4���,��`-{˨~�zY�u�������{�z��/���hn��E�6�$���(�_(54��5�Ll� �%:��o����g
 ������x�ۨ��W���׮��7���㗵$��������E��BI����䌶7{���@A��w�t�����+dcΕS�Rp��2�i����<�g2��e(��;A}}ͥd[��,�\.���Ymϡg�>������|/!F�6:���rrm�v���e3�I##�h8<olCÎ0Y&��O�K�+�� >�\Ua�HEE�wj{c��"*�@�����h�D�t�8�d��T;�R�d#�I��y�H�LBVW?�|�W�M�A��Ǔ�SI���ke_�>K�1Ĳ��D|�%mm���(�YĎ6W�X����gis������陔�ȃd?���I�W���#���dz�L�T�փ�1��A�%���n���A��G_1$Y1̫��h���M�r���+D�8bV*p԰#%D�P3�)�Ԛk�״���O_1U��͖����2E4v~}IV\;�	�a�Xr��v@���M��ߏ.Χ���W�+�%�a��f���p5:E{����ώ8FV��%�$�&(V�)VS�f�
���$�;�_&"@P�p$�nI�Q̾�m�ϖ0�q��h����z��bS�XGK��A���Nk��%q�
ze䊍T���}��9;���N.A,*�ށ����T���b��M���W�5�		�bk���:�`����.$s�6
���^�_z�ƺ'����=^��U����u����܆�?�u��+>��(�a@��q`���lo��2.g�ѓ������bsL=��`�òj�Q��Eڠ�h�) �9	�cѫ���0V�.'���|����i���#�w�T��W�'�>�E�IV��-�q��M�8Y�Dwk� ��f�u�Z�Ym�
)�D�2�t?5@ϚI@#�� k����B� �#�;�"Q(J �e;�\�\@�/�E�[����ˡ��}��Ik0|����ؔ�9���L�Q��ֶz�B{��"�[Lj��|��X9D��7���CX��d��O�`���G�FGQ���x��Umrd�{ұ����Rđ$�w�>H���P��h����3��+(z,��0�A�ʤDFv��$���BΣO%�F�솞��~���i�9&�ڣ5j8���<OLeOE9U�Y1���Ϲ!�Ž7�=��%�%L��x�M@��$�E{mV흓�����/!���S$�:�r��1�KܾԚN��d������7���N'����H-u%M�e�p��)��l��&
-�N[��(�8����u�R�o�t�O�ɒkΦ��d��d<��:���7����� ���C���D|���A�]��t�񡁲���[i�I�1'K0.��$��p�9���S�n5�?~Or}x^�;�7�#�ȱ�8��}N[�"H�P��GG֪-� ���Ct9��:���q[ҍ�����]�eZ�h�	��ΣN&˼edV;_�h�'�-?��G-�Z��j�WL��A,�pY)�}l=f�C�@?:��!0�N;��l�Vb����6�f�u������ob�`���a��N&0�Ť�9�0r��r���)0�c�b���3Z4D�)�-�����
�Z[$J��XD���j��m�dR�.�z���L#�8o�}���j��z�d�3���fGr@p.���F|�	}���O\=�%N�۠����k���c�5*l�.2G�����g�b�еۄ��w�r�TK*��Q�\��줴K]nj��Q��x@>d)J�)!9�m�T���Ў�S� ���c�5�O�2e:!��;h��!,��،�������/<y��<�'�.ްK\�6h/q�P����+���Z�o��Q+6Ѐ�-�GPN�aX�.[H�#�&�БD�f:��g�۫3�%�6>P��rɷc����h�����j:?V'<���5�������h�a49�;ΗI�h�.�K�v��2����,����l�SO�o�>@.=u��
�)0"�Y�Y�=p��j�Kj����1��8g!"$������a?gV��^z�i����6Q�¦�7޲�Qۋ�h��o��kX�迣L��N��ܽ5���Z���`e�%_i��
�c�Ъ�Zz�v�Jt�)];����؆7��O�;/�q��C6��������R��%T۵�nB֚*M�c��c�O�X[����kh�>�FA��$���A��h�=�o�ƺ�{ �옙�. A�0����n��1���n���r
�f#IBګD�Nc�R����	�l� �����m�B�ř`y]�R���b[���cؼ�-���ךa�;'� w�&��4"��qS��F��ގ�sj��"ڐTշ���'a�X-���.�kx�X�a�3��Y�&���BUm��9(�X��r����m������ћ��C ����f/��r�i�)ڋtk�/���m�bq��5��6sQtt�%�P���KlT�7�Ȓ��E�@��R��v�j'�Ժa�� ���Kp�"�2n���MG{�bh��<^�lK��L�8��a�r�	G�/=MS<QuihoQh�	Si�'�c�hofe���$o�@���As���(8��cN%�
�}�z�(�W:��ig���H��{�M��GO�����c	����s�ϕ��8j�̅�[v���N)~_bn���^��8���W����8q>g�������tu���g�ď�9��D�I�����*q�8��~�kj����~�-���M�{$�]G{�n	E�s�<Ɠ��"a���*`[�b{]N	F@_��h��)%��/�"5����(�|.1�$^�������%�z!F�Z,�� �� �h��
d�՞A�2�lH�����U�<ST��o�n�"hoBx�����������ޖ���YL�	r�^K;o��1+���(̢�1 M��/�9������_I�a��N-��_�+�x��'؂�e��n>6��R)���^m�U?\��SC�dw�w�*���~}�dnF_������{�پ�A��:�$A|k/�e?�9&L!��2`����m��h		9�OE=.i����"����Z����8P��ʖt�� �����;�\^)��>�H
|�	��u��r�&01��r)e>ڃ�Y��l�l62��9U~��߇%��\���|�Գ���`-�.&RV;h�"V��u[%��!a�ms�;�}��q�����
���d:��V	�єK��/�u�dN�p�Q���n�"�5�U���1ɓ�*�<�$W,���9����6�#�m�D�b�(c]r,��t��M;)��>5���r�6��źb ˾��&Eljd@�bJB{�,Y�C������~�e��'Z�D⬺Ԁ�>�,u�ھ�mf�ѐgw�D����n @�fd���P���"[Ñ��y�YbmNJ߲����Vy�͸X7_$�q��E�����k:F{�"h�j����a᪘m���}�#޸3�=\��"n� 7H���ȓ}!�BfR6�*lg����/�Id�JH�I�1'��
�,P9�y�iD�F]n�{e����nX�=C_��\�Rک^��s ��͘��Q�%6 #<t��X�0�2$�6h/���cx���I��!�y5�q��f
=�(E�w�R\�Jw[�� �z����OpJ\dg�ŔG�cK'�!���m"��	2����N��5<��M��V	zn���9ʜz�z�h�)K�;e㇄��Cu	&;�%��y�h-)}GR��g�"�bKs���Z
p�W��bd�
�\�m�s$x�A\�H�Mf��-�&f��o�D��P<(��}�����ͬ�J7����Z�B�7�+�qW;djC���{���dx�@{Ѱ?�"�����7��t���^hڋ�W�醑���'z�q����׻v�x!H���>�C���r1��(?�&El� �?V>d� !�q���|=��^��;y3]���#9z�x���`I$�:�xM��;QR�q��&��Y����	�ꕧbK�a�(����&QŠ~�xF=��&���b����'�zӀ�ۢ���7M%�=[U�[�]��L�����}n�}���4���w��Vw��ʾ��4{����"���㾆`�V�����Y�X+�E9J�!���d(Ek�)����s�@�z��ޗ�(H�[��9U1��2m�<Z�& ��U5����f��bO����h���G���Nƅ� ��U��|�Xd��*��L;�~��s�,�ql�����{��f3ӟw���J��:33ɶe��������^��*1r�j�<#"����w/?����M#��&�ޯ��n������U0��f�m����Y�l8	0�\��d;�4r�{�y6 �D����	�������M �I�� ,G�Ly�O45��%fQ4�g��L��"�!���`�swh�|q�L9�D�;���řϿ#�E�j[ �����b��6h�)�U�>�0{B�u����E^�(�d[q�U7ʾoz�A펂ۨۮaw�eS{ː��{W����B�&��S4hK��a�%Va�m���\\��ؾ
j��w��`>J���l�6���Ep �˪�XB�m0a%_���b�5��3�`��0Ajq���`��ĂB���)�7^&��1�y�r���.`�ez�`N:�d-L����u����vru5P�u�3@#�t���+�>�̦�[�j���s�'���\v����7�kWSΨ�T߯p�y�P��{-06Fe�5��DʆB�B�� ���i�ѓ�%�N;�^D�Ř��#�ݰ]P�	\����h�	V-��~�l@��'�*��f!������r�;567Ӣ��!���������}��O_-K77���L�2��3>��u�5d�/�?y�"�{i�)J��B�����)}�Ggwz}�	<��JF����ޭ���E�~��2A�g꩸�z#q�UWsQI���y�������)V_���Kz��RQF{~w!ݷ������U%E��H#�d���5IN��\�l���o����v9"���j�9AJ��K�{^Jrd|�5M���V�8K�<�W+z�^�)vN��km�������7GG{a�lwc�DF ��~yŬ���������kZq�n�Kh�^؇<f+�ܺ����`�}����9it��Pu���8���/����ҭ�b[�[�cu"���W����bv�+-g���-h���;+$�2DV�h/0�P�����NXǂ�����Z?����@o������&F��A�VyiI0F�ӵr�^nR$�A��P�u�~S�Qb��t�]�+҂`�qCH��>�4��e�)a� ��A�`�.��`�PX�ơES��;�[���b�I����nWy�c�@����ab,Dȑ0s��y�>@�,;]���= ��?�Fi[>���F�n��0����Sg�m�VHl�_4�"X��@v�Jkj$�OkΣ}�QDuL��+}�:�L�Dy��i�+��j���(���.�vg��A�ZW� +��J���"��J�?9��Lw���/R��O�,O�ixzu�F�&�]L�uL{�����7�e�\�=E��)��!?;ۋ��VS��z�t���ȏϤO?{��w�eU[�0���W2��_t9���;��Ҷ�7�N&F��NwVzic0�!1�f�m&J$�N���'S��%��a�a�h*VgP;��?
)�ڠ��w�s��8�f�����!���JҊ�!����V����3~u��]D�H���?[�K-�:1��b]"�����Ĝ�a��(f&JϪ���]�t���b���� �]��H4�D��k�N���(gK,	�5�g���Wм�hİ�c�Aإ�'!������pC}�u��бl�z?|KK�a�uG3��rN1�ublbt�V����|��H��n<DaB��O����O�'�GSl�Z�n�ў����y1�ߖH�V�,��1a��D�~�X������F��\���J� �L,��AcM�/�i����e�אo��kK�3[�50Y���˶`I��ӧ��6��}^��?b$6��f��L���䑹��w�܋����"!��O'K�bj~�~*�Ui{�Uu�����z��\��f�؆� ���-�K*�c��'_8@��W�L���=�uu��0f1�
�����O?I�l:���{�L�ܱB
~�{�7�rݍ�����;�g�fb�zIU�(��(n;��D��Q�.��M���Ɯ2�̇S$��1&����;.S�{���bW���;_����aګ� �M-uRL�"�A��ݪ9��������IX�O�#ţŮ)$�t��S	����jw�bl3�>*�EbD��a��ѭL;�G��f��a�=7�9����ߑz�&ݦh�-�x���R���{�f��2��"�<-,��V,��݇j*wa��fv�?���,��K�nEA���ʰ8��،Ee�g�祿pGN�tF�����٤q�ވ���0��7��a�?f瑣�D�9M�E�ϖHNT���XJ9#�Rc�"�\k(�#'-��iNrz}7��A{[���wn'u�b7���gXƙ'312g Sp��q�8�3?d�ɤ�Y����;$(�����7AH>p i]W	�ؠ���R�$��@�yL��T��DI�_� ��ʦ�k� ���70�Ⱦrd����V+"�?c��Of����D�#��'�������*��ׇhؿ>���g���(�����$�	�}Z�`���ڻϒ*A�%a���n�QЇ��Ĩ���i��,��i&s�<�����"�jU�s��zAr��'_���.���߲�ZE�~4{s� 7y{A���j:d�jM$��E�yl�(7���3TT<��/��j*$0+��Fv�����[��к������ub�����Ĩ;��0����r/s�]Y���P��$j@{�����K�{�u	��4�6���B*��c�Hb6���'h/�2$�e����o�ꗧR���P�駰���N��(̺�������şx���1�31��Q��@��(����9�n&J��E��u�w�bm)Y���v���,��x� t~ON�&��y�쮕�q@&A��z�>{��3�01f21��GbDY�D��9��\�i�ݿt���&'L0{p �۫�U��ꛤ����h	�Xȳ�>6m=lR[~ ��p>�"t'�����k����������/�tc~N���t������1fb�����K>dU���h �!����ȡ>Muԓ�q�E�H��ĲB��Ta�-��L�S_7�	��mшt	G���J2ڸF����b|�Z��j/���0��	Da�u/��~E�^�.�'��]�K��SU`�Q�ho��mVb㱽�^\t�Ԙ�%������Xq�ؗ�3ݒ�V���8�e{�n1�����~��0��5�;��g�gSO=��]�n���U�'Hem�N4�D���L��w�����e�H� LMTib�#*Sq&�|����_Q$r_sv��&~��RfED�Y�Ʉߕ�4��K�ʽ�y�J�T�D&���0�R
��v�יACP���v$���)�h��Y���w���=L���2���iV�E�?D�&��J���������7&�=	h�|<�?�dQ���Ȋ&7�ӈt�(�է������)�������纫�/EP�����]!&J�D���su�O����4�aP@{�(��% B��f!��SY��@{�o�yn���n��c����2�fD=���^�+X��CG�ŴRd%��=��`KC�Al�b�O�B��~"�T|�)5��������^����D�G#�o6��d����yz�d�����=sUj�k��<�Tjz�~Fjn ��A�#����]#E1�1�ck0��/=�IP(�ml/D��i�X� �ɥ�$�l���.v�<�42�g��uC ��;��N��=���0��h�"R��Px�BR���Z5�05�{��/F���g��0B ��b��x^z����?_)c�bE"�Pd�'c{�(���A�)����/�DY�u�����a�"���f\�+o���G��G�Kx�J��{�5ٚp��?%u�\z�-+d��_�{�Q�W���'�ȭk��㖣E� ��g�҃��	�M��)�\H�}1V��}�����b�i#�?x��	Jٶ��+!�,�5�Lcb�g�����|�$�?�/v�x8){���Z��l�.A0���ˬ�iV6�����Z��/%��^d5�=���U�uW���bZ�|ƍwJ0����W���� 5H{��b�,�_�
x�'{���{���B[����`#\e���84i����U�`��oO*�#f v�n٠%�4� !f8H��*:#�@��8��`��b�cb�k��P��3I *�/�ޚsOd	q�dr�y��f-�+5WV��P���x�n�Ò�u_�[��M��3��^YZ�!���-���*�Z�֣��i�6��Ff�F��( F���S���a�LՀM�-����7�)ɔ���dӸx�N�;D�.Fu�i5��)�^4c�1�`%�#�v�@��̊QsφD9	��DyDw�>	�Qb3g��K�B'��S�4��a���^G�;�����p<�h�h�Ѣz�+��qCf�h/m�Q�׉�sJ�F��� ��G��]$Fb��hU��*p�����~�����n� ��Z]����m�@�c�Y|����b��EL�1:h-�4�t�C#���Q��X��7��^�X-�?+3�
�Z�t��/h�QF��L�L��
\��*y�g��ĸ��OC�� ��R��.�s����^�ɾ��_\H_��n^N�_, ��A���i7�J��P���p�����D��D�� ��c�4OD1�:�t7sF#܋� '�����P�B�Ba5����S��E���sH��E4��Ǩ�bYؿ0��؞ʌql]�������o!����y�.Z�eJA!�S�F�꫇�( �8���f����b K|UO���\��;G2R2AfA1���s$G��_.�

��bQ\�~�5�p�,&�v���æH�������Κ�2e���ȋ�&�'�kU�����Z���D���IL���)X_�?HK���aN�Ŝ��Cb������DǢJDl�:*>H�At��#��|v�uG3�<����7�nb{GS���J��ĵ��۬�"�-b��m�D���Ɲ[V��)��X�0!^!sA�8I�۪�B�	L��
]�R{��bLfb���Ho��b *3�r������xåTV�o?P��l���+!���Pc�1�43�G<�ޢ�{�v0��ڷXb{~�+��ᰘ��ia��Y�݈�_E��C�"�q�B d%T���]�M�qL�?1Q��Ru��Ę�f�;���z���MO�g.,"�GoS����%C)Vԗ�i�U�'/�a���ex+�r&J�#}�b{����Uī�5���p�.3Γv̌-jm#���AΓΐm����/�^���ۛ@�1L���()���Q� ƏҬ�Gv��zJ4=���W���t"ȷ�G&�j������'x*��-D��s�ul�-�e�RzV>���A@�Y5�4�eA�Av�KG�����nK��[��l�L�EsY\Q�Oϗ��?�X"�(#�R�KD1�rY�V�Gc/���6cJE�[j�v�!�{�5z��=���5%[(t-6�`)#�5ڋM���4v�	�ͬ�d��Ę�b�e�>���_<-ʊg̤�ɼq��2F����ϕRq茔͎���$V�TѰ�z��K"��z	b�ĸ��ak��b�!�jNe��g���ͭ��;t��T~�,sLj��b7��SX�����U�c{Qp�o�Ш�ߥ��'Һ�_�K&��,���3��ch���T�9Z� ��3K2zY���B��٣���)���( �	n+�l�����E\C{�R���Ȋ)�D�'����({�|kQ�U��Xi�E�;�`�k%�ߵHQ�u+��ki��OS���a���XW��)#��FM8���A�w�@���� ���D��(�T�Dy��r+����b��n���>27�21Z:K�ݥ�y�I�������n�9�dc������A[ (h�uۤLE����9�)�7x��4��_RP/NlF(�b1��v����~ 7{&�gQ�D�l�"Q@�ә�3g�1�f��b�%%�%�E�޼�j�z�R@�Q!���$��!������*�%�P�l���j��"F�S-D髋/l[�j{4,@�?ɰ��L�6�Xb��o�,�.5����RF�Kz�.�!$���e�\�R�jI��\Gt��D	0Q�:�=�)�8��qCeb�� �7E3BJ�l@jc؂���v��KJ���dePCs�����PV���_|�<�}UK������Q�$�����8;�NW�|2��obh�?�))x5��/��M�h���p������^As�K;6.�`�''��N*>���m&eJ��+f�{��|x�i��
F��R(�3��,]�Ĉ�@�N@�	$�Q����D� ��%��(��5c��O�޲-d���#7ÅdZ�,�V}Ku�����~O������_��[�%��r_�,������#taA:]��(RS+����ZAFk�������p�����є9���A2ڛ�F���/�D����O1%�'��-U{Ki��h�%ג��H4�e��J�)Z�p�����tߧ��U����ƻn�Pݪ2��N������U���e��b*9XC{U�s�����#��Gl֜�S�ьY��9-h��1�׏���7R6(�Cv�� ������5vZ����ܴ�&M:I��r�VҢ)z���V���LFo35��/*��~*���y�7��r��^i�7�\\A�m����K(�n5?6�ʆ��Sx�ץ74���pI`�jRv��oP���B�����DՃ,��:��k&�"��߀�b�Å��?߈�Ϳ���x�ޯ�h�<2�MYw=JP��)��lj���lAR�ץ��u�Xjz|���R�!S��)8���9�G�cO"��^C{U�æ�?�����j	E>�-h�Ί�--�$��D.Y�7k	�u��%� ;[G{%����u�8�쀌�H���1����'�>|���hb�t�?,C`��u�H��n��]d�i�����&�\�mQ�Ί8,���tK3M6rg��f��l��q����]z�������hozF>e �ݹM���
o>[���λ��Ƈ�n�`���Ϊ�hY���I��K�SA�l�@a4e;�i�Hj�odr�KFC�6���+�W ����5�I~�%�})���;w��d�ُ+V�������q_p����%��fy�F+ʩ��s�#P�(p�n	��MP�?��#]jG�4J��y�'��~�U�K|�uw�d�:��;��x�ukiϐ�G
�_�n~���p�d>v֛���+K�IV�24��a��;T3q'mX�5��L7�Lӵgjh�q3hܨ#����eA�@{Qa��D�%��R�j��>�$[+Z�C Mn؈���[�}�5�7҈7̼%�[u�����BɄ� C|r���K�,)&H1sãr��A'�ł�^#Ż�,X��k��z:��ǩπ�q�W�T��M�̣Q���%���[(�件�Zמҕz��I��ȶM���_"�)3'��������l����=Nڻ퐡R����T�{[���@�h/ʙbaeȕ7Ұ.��U;сBVkVP�̟	���D+���3�b!'�m�ᬀ�{��Q����k~�qB�* �0V��6|❌��	� ����Rj��ް���P<ȺS�7�iU_Y
��I����}{)�o���U���S�oj�u�T�Tf���6KW��?�*����dj��7���o=��+�fk�B�F���������o���$:q\	����*-����i�����t���B�qR3r���h�A����V�2ܒ����uiz�fQ$�%8b��~Ţ��\|o�.q]d�+��8�M�a#%������2p09�=Y�J��?5=e��@:�{�X]iHz���(�����Fq��-)�V�Pg
���<��wp�G-��J�߽���r�KA�3��a�����k	��U���?.���2A���ް�G� U	P���#kj�����I�|^���em�A"���n7�v�L~W����R��@{��j��䀴BL��'L��H�~uy��ͪ��D�>0��b%���RP���AbB#�����xx�Z�ab�E��[�V���T]@�]��噘����q��3���3�E#��n�k/�|�I/H�n�!lanС�KKU�j�ˢ)_,���5�~��ɨb�UŞ�<G�{��wu9�}�w+�@XO��Ȓ1�p�_"s�J;�<��M<��J�sN~+����D��oJ�;& �\h�B�FKXkd�v!*�Wz�	ګZ�J�yh/;�;��4%������
��8��Ye�=b<͘5W+#��Ɂe��������Eו��јC�c���\s�ށER�ߩ�n!8�>O�vZ7`b������S	�A	l���R�-���#0L��H������qXs�n 2B���<���R޷^��?�'D��F����饗����y�O$���֫��	"cS7�5�~�w9<z�F����S�'WJ���^�l^�a3����jbƎ�>�5�WA�Ij�HHd�U����E����0�;`�Illn�T�	.�/�W���4�)K#I�s>ƠpF���� ��̭��Z�>��	g�(�OOI|��'B`�
�Y�utU}ߛ���;[�HB`Gf��a�CM*�����K&�2F4^�HG{�yb�)DF�!3+�̻�5�j�?�L�Έ�:�/����N���>�G��DZ�s�h0���T/yT{ᙔq�L��(����9�g�݌҄��Ҽx�]|	�5�kdr�9��ЊY�����6��'�Ɛˆ���v�&/8D�a,���t>5�q���6��gk��שZk�u7�f{�����y���*m�����b�\�i�YS/���9�`�I�̻���e=})/���!��K�� �E�I/<y���;Q>~�d�p�C�r�������&��Q����n��D(�O���Μ�Z' W����7Ȕ�G��b���i�u��7b��q&J9+���C�@)���}�m���� w+��v�j2�� �`���5[Z�8��f��ꥱO;���ܟ�Ϛ.Vć}S9�>�'[�����)TR@
�����o}M�=Uz^0�oGh|�v�E��lb籣
_բ#����Y�$��5ڋ�%�b���{cװ��L���H2d �%� ���D3d|F)��H�ٰ)F���\�o[^��`pA�CG�C駀j&���,R�"J��"h/$�¹Z���U�Ǝ(��w���b�m�2g[�ETE����|1�br�Rz"
���Xw�%�=��JN���4o�*[-�v�����R�X��-B].H�����O"ˠc)�PF;�+(ĺ؞ʗ�HG
Pb������S�*+V�%O����z��#���c�a��_�Z"P��J+�A�B�1��B���+�(�8�Q�R���{"�G*p�^�>]}��}`v�������S�h�6v0�8%�U�7�����7L�/o=^+��,o6ۙ�-Q;�)T5o7����>�8
k~u�V�v?�V��i?����.|��q�8]�IEQ�Jp��M�����-�D�:��I�������`����(�o��>]j��/@�S����>}�o�nz�ˈ1�Y?0�~/l�9�����f��c�؟q}";�k9_�f�|��װ�.�����L�E�O$�k/r�w<�"������$�[��F�ؘr�I{/�<�d�v��,/Y!Z�ݕ��(:t�^\�=X�Y��_C��ְ���\( �G����4/����\.��e�����Ֆ.��8�t
�~W���8֐0�?�pR_zZ��'re=G�I�h/�����Tկ@�^ㆠ.v �$:�X����i��f��8���h8H��
~����v��(˥�=!u8�I<�D�H��U˨���o,�u���I��H���MiO�L�Q��
�fQ���I�zK01� ~7
K�O����o`��5��Ţ�~Nƅ ��y ��)������K��#@��YM�SI7��B�{Ļ�"l�[ل�0J�[�� I!z#|��$���ӦO�����>�$�K��(�����iDk�O���Wҏ��a,�@��}�aO��0w�ך#�����D��E{YL�h�.���)�m�521�\���᫷�f���#"�Ac�e����S}�29�޷��u�(C�2�i�H$ r2�NI/EI�<w���8uuk(��l�_�s�EYQX���@����jؑ�����kh��(%��z�Ԡ�!��V�8WR�^A���>y���t��z���YO���T�=�K�C:$�rLJ�e�|�� t&��'���r�qSE5�_�XGdy�+�)$RBW�+��1���5Qtq��n��:S��^�c�b��ؠY]x���d��a�W,�[�� %ak���h��ﱓ-����tk8��������F���R���ąx&T,�?� 88n���3���[�΍J3F&Sm#��Y�4`j;>�&���ġ���i�h2�iAr��4�P���Slg"�;�hXlKL���^��[����������c���XA-u,V!���dg���(1	�@U`W�֓P�E�'�z���^�q�菁àa;ofm��2c��x�dqh�r��ŦG������^DC<�T�u1b�;���bTD;�0�6�~i؛�K�����f�_�:c���8���K�9
�֮ ں�2�Q�#~���?�ܲY�!fsṅ�x<�m�^��-޺[�0>�t6�>fn |�.ab�D��m	h/���-� <���`Q� 0,-Q}�[hVJ�Y�h"���N�/��:�X�׫ڶ����4���`	����R��_�A��Z�n�eA{���9�n���<ـ���
����\�ld�i[>�?:{�I��b|�e��ޒ� ��iKe� _��0z)�'k/'y BJ��R�]X���Z,J�CF�Av$�8�՗/`E�G� El��I�?J�c����kl�<��G2A^2��r�-X%� %ڋ/&~�T��Y��G"�[]�U��6�YZ�?sFp�Dr_�[�`���lfV���/���n�/���#O ���h}G�T�V�kWhK��d��̙M���h+�z"7/�Wo����l�".K����=�4b�&���`c�8h�� �������7�qQ[C.~��uN�9����rP0�5w�#:hL��P) U�edb؀��y�>����|�*v-�(M@{���;�e���H���t��
;�If�t��#�V�`�m7ŋ�e�/���+6Q~F:��n
2!{+�!�LX�?��CVx�4��	�IѠ����um�������Y�x�f*�ʤ��t�5�߹��Ȅr%�=~��:M�x��]5��2 �^�g;�;� ̊�)l��Kt ��p�N
m�(N_�i��TUUQC%;>��a.ߪ�!Q[:��\D�ۧM�e=�ۻ��B,�3Ρ���4���i�ІhvQI��g3���69�Dol��&ې�F��Qh�z���O�ڒɁ����)��)\RB�!�w�]�]VFM�x�|sfu3�
ƐYJ �8ī�ָW ��� qDt�����U���d����u�{����FR�u$e�Tj��X5�)͞F��^��
5��lK���4���B^E�n��+��-o�I>�V���ʠ�c���G�A�g�����[���*�࠴�<�Dr�|������U�]a'2c�+M�_q-��Ss�UR��0�$o������z�vn])��M:x�hż���|�r�M�V��|�����)qx��5�}<�'��p������[Ѳo���Л�"�BA?m]����m�Sqe��6���xZ�K�7���_1�Ɂm���������%&��7��h��O��+o"��/�#�eM�o�B �5+(��MJ��}맷�Y�P䟳��?k��D��4�J����*(H+���'�{���T�eu�b���i�sΛ����+������A���Q<�����\����7�u~zc�<,�f�k�U��v2\�����kWhA�Xw����̪�?��[�;P۹{@���<�����tu���\�%��'��_����M���=9�!#L�Ŧh�����=۩�[Kӏ�pZ�L�H�|�FS&�"/"tEG*��)��j6]��]mlSe~����ʺ�cC ��}d�2�	"1$",$��E��	�hX�%� �?�EuL�&#sf�}�)h"$�#�97�n�-�]��޶�s��ֵ��x����=�=����9��D5��U�й�F��惰s�j>��r�3-�%e�N߮m�DXT�[ޞ*����1̴.���W �R�>���<��1�3���I6s=k"q��;H
��ywV���I�`*�d�L��+�g�6kBd.�l���7(yt+<{_C��S���ܫ�^��g���a�� 5�	j����N�ܛI�MgGϻ�[�߆����S���=�e�v��!�č�ptO����
��	�2�H��Z��~�p=?-I3HO��L E�c\!�m��h��/�n��Ȃ�q"e���l"�ڑ7�C1��jk�w��Warb���m�#�5���*�-�S��
�����+a�u����F��^ý�����S��l<�JKM�2^�U��IZ�j7�>2�7 #E?^B`Wb�Lt���� �$�����Km��EJ#�`p/��밷�O{x$�ݚ!P�n�-��`:�bf���_�[��"9�W�����]p:��e0�F��~!%��2Q)"���8���H�y!�Tp�����l6���Wj*u�]�dr3���8�W�Q^R���.��X߄��=��w>��� �~����6��D8z�d���{��аI
�3���n�#�d%V�B��$�tm64��Z��О�j!��-��������0�/��u�t��yT��$��b�V�!\~��B5�ll�cO�6��%�89�B�C����O�k�r
��'jT�l��o�Ů�\P���I���O��Q���?��G0�R8bF����a;| �������^�!���OVF}�#�3]_�r�u�͐�Ԧ0=2%npae�a����;ڸ�	���$�ىt����x~�š�P���mQ��"'� Wx�P��#�?6';O&�<-��z���EH�l��h8�J�*p��,B�7u9��X]�����s�8��3W�!����A��X��UB^�h�mu����}�a��s���9��6��:i�����&#%�o��l��n��\��X*c!�� {�~�Tw{���h4�2�sW̓��:W�[��"&�ي�/7�z�.L+I��KlN8C79v�S�[���:�ǑRb�=�����O���˅i��$V}�um��̰�(���,�\�*�[�h��Q�����(����Nz�Ø���8j���l.b�C�zE@��gޱ�� �Uŕx\��    IEND�B`�PK   ��Xbj.�  B  /   images/fe3f9adc-aa37-4826-b52c-f1f60efd89e3.png�XWS۶�"�@(J<���P�s�)҂ r(:��r@�P�%(
����@�����D���P����y�����	/cd���k��k��%��Ԑ�G�  >��������'8����/�n�L�@5������q� X�#��2H �i����<ID���۴k<�c}��T�ΰk�6˱K�it�����f&����sT�B���7�q�F������b�f��+]st�9��s2,�a��fB�G�]dje2����Z�\T���^��~u6`��B��I�k�nm7Wr Z�?��ɱ䝞m9���q�+8������p[_�5Nj�w���A�C��D�3��z�ғg�c^��Ҋ����Z�2W���k����Q�|2���JWA)A���1����F@5���x����1S>Zc�E:^5���69Ҭ1|��i]�H��4i~��FaF'"�n�Db�Db�]y���>R��eS� X��-V"�D����Dƭ�W��F��R����i���RLyy�Z�
8��H�~1ԙ(��iG�C �i��2�a��~�x�Y<�~�f{P�:Y9M&|�CE����|v1��:پ��YxIfҚF�R:��҅��:���j��������8]�(���CD+Z�U�9����}���\��&=4a�S�"c0J�dŪu�f��j���W����^J�>Hm	6]��P,���'6�P:�r�j�Ɖ�1Ey�%;a�B�e��D��a�D>�'"B���?�F�8��,U �z����ٵ�Ӛ&L��_n�����8_D���e�}t����w���E�w�W�*e�J^��z���}�W�n�-�mY�mA�=�Q���b5\��'�ݡG�HF�k�����q�V:B0�K�-��q���Zؑ �G�v���?_n��1���
��z���Q�NW�+%~4P0քK��u3�l��+>�P/�3�Y/�9���R�Z�)��H�b��s��k�-���.ြ<�yԆ�O��X�d�6��|�o;�mn�ލ������V��v���2��P�D�Gd��;�nq�w�ܸ�pUoBE�3e$�����+_��'=�^k."(�.��dG,kiWSw~&��#�_�Q�0�Cd7�9���d�?EDB{�QWO�gkJ$چ`N��9x���+�E4v��\�io�XZ�c]�2�Kb'���K�j'���r�ݿ�5�_����x[��A� �D�T�)Uy#�����ݾ��d�Pr�O������U�e�.ck�F�"7H VG�q��i���c�'D��H������8����N�;�~a��׫�,6�)8�5����*�_�e����,p�aH��W1�+z5�{-�K��ìb*��g�����t"1����tʏ��,��XH��z���|��RAM
�H:���k[{��o��˪D�#��*�������D���f����>8��K˦}���rH�3	��IC� #��8�P�o�X������P��l'�����Ge-�/����2}8[�q�Yq8Ƣя:OiH�����/�#�
i�*�w�@3#kB;���o��Q_Jx�3t���7w�:�惊*����{����ZL�~�P�~!u{���KW���kۯ�JW�Vq��|[���v�WC�)�
��9<��`�g��dy9�������:�/��Z$�����v׊w�����礚\��ihڷ'}LKR���R7����;����&�+-�uO�sv�wf�g׌�0�L̒������*��X �Ƽ'�.�d�m����Ə�m�6�]O��R�*��B*�L��B�M�ej�Yl�flyi"�A�?�>)�;Q��_�|Te��/C�ʠ�a����m���ð��6I{Ú�M�&�Y���DAl��GmU���t��KZt��|��
���ETPN����e[�3�*I�Y���]��7�|!��i���	I7bE�&��]с�1�@�޹��w���o:��!����
@~�˛�9�5�X9揮�����Mi 4�_nPSW�8S���d� .��ũ�ՙ^c{ ��TA��� �W���pU��*E-�7�Za{�o8x �补N Խ�w>+�Р �U��2�����л%�/g�
�����_��!�2_����|�]��b�d�>+�o�*���l՚"�$9�����e3fM7��{��)G������t`8�>�v����^p-3
;P��!����c^Ε��y�S��Σ��F9�陜�����k0�^��3���皇hd6�`�U�� PO�����]��3�9��B���=�C�L��o�X�썫 >�� ՠ�������%��2�O�0�#e��(6��O�, ��|#Du�qq���v���d#������=����y\sh���q�}$��_�ć�]��Y2��8�.���E��U���eg#B�w�_D�kH��0f���$��
m��R�Q�6J%�h�u��@��n=�x�U�r���k�-�b]-�<��7Yω�z�s����+�������ea(�ރm/3irƭ���NXV�Z���E���i�O���I�eC��U��^�sn�5\�7a9����)8���,�a�=�O�S�����6:6�-))�`��V�F�c���b�$V9ZvG)�����>����.���G�����놜k��Y�&��y�t��(8�v����Ҭ��
���eF,�7<��u�ָ\�.E��5�Qm]s���%pEڜ��3����O��rL�`t��h�o��I�1;'+;Zh�8D��U������ӊ,���3#y,�iz��~������Z�Nyg-��4���`ߴ�y8��J�[�f�L_�Lw2�G���<�.j��>q7 ��M'��w�&}����@��{HB����U�{8��>P��!�������U�E�-Ҭ"����g0 �cC��JO��0gO�xϑBD�]������fwA���n���?P2^me�h��R_S�y$Z)�sͳ���'n=�G�Db ��H��y����B�pN-��e=��~C�q~|<}����Y���2�wy!Xacq�:��'����Zy�j���.4�3���c\޶Z��a����]R�G���|��K]Z�������ܡ��=�����d�`�eʌ�S��#T���{+�Zd��)'��%�~&4��%c�(�l�]�:�yN�PD�ۢ�Ão7�@�d�+��7�����d&������=��F��h.hR�ˊ�6JO�aZ�����K)����H?GRS"KE��O��X�R��(��J���(�)�ޠ|C��E+�=��0��f�~勏��üg�Ímj���(r�o��KE���U�����_{�hs���������P���"*��y�Q�q��Z��qH|=���U�O^����p2�ƪ�W��,&�`_�Z��zׇ����*m6H��<�.#�ڎQ�	���%�l�^vchs��_�cd��G?�x�.���c<�ͥ���>f�Put��\�U�6�ypo�[l�^MhX�P��#ټ�4ʦ���ٶ�7nEn��)����O�3M��l.��R��0o�E�0��1!Bi���ї��:���~�{�4����D�OJ��7i����.�`�H22�t�[�J�Y1�\KGa�2}��@���~ݡ�\�YȲ:Q4Ǣ���a<�#�נ�i�^��%���S�����	��!-߀oO`�mX^�إ�=4c�xV��-l�����Ɵ�-�ͯY�m�:�nLɭ��j~�Y]$�w�7|NU�(y�I�߿�!?/m��x�i+O8�<��	����oJ�ݳ����B�
��f��tBڴ�f	331�t��8����K�1�p�j��(B^�&�1Y<�C��(��[��lW8�����;k�ʻ��T�c�O��;:��ɰWJ�h����~�0��bcg��z��G� Z�3�ųerC���+	�i�_vv�T�g#��V�.W����؛D�BV���#O���@+mАS8��&��J����P)���L"��m�/u�2�pW��X�.�L'FX���e%%�����Mzf)E7�q�7�c�<}$�7��`:wP�}-,�1DLE��T^�J�3�!�kIׁ�>���̣�J��(�Pn�&Rx̤�1%�'#�$�p�%�Կ���w(�]��{T�{ ��ӡ!�G-)��&�J��$��4{�ɳ�����t�'�6[�G7�al3]�m�|��	���CZu��	�-�k&�:3��2��G�o7�ܵ�������X����]��α�wVz����ܴ�-<b���)Bkisg��m�8����w�����d�.jf�a�"R/��K$(����I�Y�}Z�׋��<acy7��2H��+�]'S�y˓�z��	�6�V��dq���tu����ҺO�������֝��]����n%�eF�����f��r�f��#9ͭ�N.Uz�}��$l%�x��֩�3$����s��V�{�!�des���������,:�(�(O�/k��D�nd�I���J�-t˦����(D���k�e~����Աl�i3��B2�<�$)�?���t u !�'���vG���d��;�W�ePj���2���I[Yk=�����
p$����ܩl�}��Ix��_L��ڒ ��}���g}TM���L|�Rd{���ѭa�
���PT�Is��BR��m�M��3�����xr��U�Nh�tOG
ʴZ��/�%<����չj� �Q�y��gg��Z�3,0up����-V����G�k�� 9&�R� ��5w)J��I@�/*�
M��uuu_��ۨ=������/��mv�K1 : `n��l�'�Y_6`�k��0��~�n^'J�?r(l�����@��բ�6Py8��
��Q�WS�.��)w�uϲ���cAq�כ�g�b9�ŤY��b'��[��Gd)!�t�bQP/}�n,�k N���+�����2�`2 ���lV�A!`"fE�kk��>�&�ױ+ ,/�V�A� `gSa���`$��?�k��p�nDҤ�˂��c�����ǉ���dk0fč����:���Z^�T:F�:O%mZ��G�,3���.�̙ͭx��	��!<�y��� ��~t,sy2K-�65�@�͂�A; ��r��
�;� ��#���ǵ]��U��Rʡ���A���(P�}~m_ K
������f�N ��T�� 5'����vlY�4��Av�Fז�ѿ�.J6���q��A����O
_�s�Т,�YC׷��AM��d��7 ��^n��,���>�+������N�,\p��̃���ʬ1a���H�oJ&�ѱ,��K�2J������y2������`�v@���} ?F�M�+�p��PK   |��X��pw�  �     jsons/user_defined.json��n�6�_��;3%Rs����mm�$�
AA�T*̑\�nP}��̞i�-ˎe�J�vr�H�t���wH�w�ř���Y��x�M�fF;c�)�4���{D�rW����/���z�ܔi9�{��ss���]�sY�ʹ;��7��
9�����LH8���'��*R\n���R�l��as��U<vd�K��K���'q�s����"H"㩣Yvc���kR��q"��;�4{�%�s��:\��"K?.�|�R_̋�>k_�*w.����L�P^�S{�P�VJ�3�����dz�6��--O2�!/lI��X�p�26�6�|�eX(�#�kf+��j�.[�N�r6��O�iY����y~W���G.W]�6�$㩱��̊|f�yZw����|Q}n�����Tu퓜.�E�[U��~��_����β��v����|\�Eծ�s�d��evc���=���\k���]�)�2���~�fO�eϫ����[^���,ϖ�^�ku�>�:�v�u���7�׋����d�\f���ķbc>�U���l�L�+a�6�5��-7�d1��ϩzLDQ����yf�����U��7���Brj��T̲���p8� G�#��p8� G�#<������/���<ˌj�����̵G(�y��/�ӄ)�#BʈPɅ�4�Բ��v@_u�A^�(vEI$��0C�C[!"�Q��b6��b����$��O�C"]7$~��&ҾX?�Sq����;�5�-༆�6��!���1�~O����������t�{-q���������mǻ[R��w��\��!\`�$f��A��p8֔�;c�5%� �\�p.�� �\�p.����q�̍��27��4�p1�ş?-�ћ"�JU��x��d�U��ѥeh_I曈$B�Ę��ؑ)��BΔj�e�1ա�	D��1�D�^5�I)廡�����+<�����?
"J1|5�bL����������a[�n�O�ϯ'�6���蟿�xq���lSBT���puzک�z��Z?<��w������C�^�|�#�k�C�{�=҄=�ou�]y�S>���Cm{q�k����_����W//κ����#Q�*���ew	}��xB����	^����mz���3�����6�C�wv˷�m�v�I�-߆��
ׄw˷�ݴ�@k��n�6���Pc�t�&m�����I�ozmp���J��ƶ�:.���`;x`?��;^��3��.ߞZG6�rU|3��e[��ɋ+��
X�v�r��;��f�Wi�V+����V�2[$R��)�
_Oc���{�q;oue�R������,��L������|��s,ϱ<�W��p8� G�#��/��^��?"ٍ�R[Hm!���R[R[Hm!���R[?&��E*�X��p.�� �\�p.�� ��{r��u�3$�~�e���H�����ܕZ�r?��\0�17��P�-�������Tj�Q��H����ҷE^@b�)��$pM�#a�o�"h��鸠��t��`x�����og8�Ӊ��o<\ԁ:P�ߠs@�1�\�p.�� �\�p.�� �9IdG��eG@�uߛ:l΀��9�>yl��#��2lΰ���؜�<6g��؜{��L���(�Ş�p8� G�#��p8��M�p��PK
   }��X�,�KƘ  j�	                  cirkitFile.jsonPK
   ��X1	���  t  /             �  images/4a240ba9-1e57-4d57-96d9-193d1ad0babb.pngPK
   *��X�����   �!  /             �  images/4b131f3d-bb43-41b7-a007-3fb3641e8d39.pngPK
   *��Xj���(  *  /             -�  images/6c8b06c1-8935-4e1c-b7d7-4989f9141afd.pngPK
   |��Xd��  �   /             T�  images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   |��X	��#u } /             j images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   |��X#�@�9� �( /             ڑ images/bb1d7dd6-69b0-4e8d-a72d-bbaa9fc3070c.pngPK
   |��X�ĩ�xa  na  /             `� images/c9c0af01-d4ea-463a-b9af-0ddeafc58269.pngPK
   ��Xbj.�  B  /             %� images/fe3f9adc-aa37-4826-b52c-f1f60efd89e3.pngPK
   |��X��pw�  �               �� jsons/user_defined.jsonPK    
 
 j  �   